module tt_ihp_wrapper (iovdd,
    iovss,
    vgnd,
    vdpwr,
    pad_raw);
 inout iovdd;
 inout iovss;
 inout vgnd;
 inout vdpwr;
 inout [49:0] pad_raw;

 wire \gpio[0].gpio_I.pad_ana ;
 wire \gpio[0].gpio_I.pad_in ;
 wire \gpio[0].gpio_I.pad_oe ;
 wire \gpio[10].gpio_I.pad_ana ;
 wire \gpio[10].gpio_I.pad_in ;
 wire \gpio[10].gpio_I.pad_out ;
 wire \gpio[11].gpio_I.pad_ana ;
 wire \gpio[11].gpio_I.pad_in ;
 wire \gpio[11].gpio_I.pad_out ;
 wire \gpio[12].gpio_I.pad_ana ;
 wire \gpio[12].gpio_I.pad_in ;
 wire \gpio[12].gpio_I.pad_out ;
 wire \gpio[13].gpio_I.pad_ana ;
 wire \gpio[13].gpio_I.pad_in ;
 wire \gpio[13].gpio_I.pad_out ;
 wire \gpio[14].gpio_I.pad_ana ;
 wire \gpio[14].gpio_I.pad_in ;
 wire \gpio[14].gpio_I.pad_out ;
 wire \gpio[15].gpio_I.pad_ana ;
 wire \gpio[15].gpio_I.pad_in ;
 wire \gpio[15].gpio_I.pad_out ;
 wire \gpio[18].gpio_I.pad_ana ;
 wire \gpio[18].gpio_I.pad_in ;
 wire \gpio[18].gpio_I.pad_oe ;
 wire \gpio[19].gpio_I.pad_ana ;
 wire \gpio[19].gpio_I.pad_in ;
 wire \gpio[1].gpio_I.pad_ana ;
 wire \gpio[1].gpio_I.pad_in ;
 wire \gpio[20].gpio_I.pad_ana ;
 wire \gpio[20].gpio_I.pad_in ;
 wire \gpio[21].gpio_I.pad_ana ;
 wire \gpio[21].gpio_I.pad_in ;
 wire \gpio[24].gpio_I.pad_ana ;
 wire \gpio[24].gpio_I.pad_in ;
 wire \gpio[25].gpio_I.pad_ana ;
 wire \gpio[25].gpio_I.pad_in ;
 wire \gpio[26].gpio_I.pad_ana ;
 wire \gpio[26].gpio_I.pad_in ;
 wire \gpio[27].gpio_I.pad_ana ;
 wire \gpio[27].gpio_I.pad_in ;
 wire \gpio[2].gpio_I.pad_ana ;
 wire \gpio[2].gpio_I.pad_in ;
 wire \gpio[32].gpio_I.pad_ana ;
 wire \gpio[32].gpio_I.pad_in ;
 wire \gpio[32].gpio_I.pad_oe ;
 wire \gpio[32].gpio_I.pad_out ;
 wire \gpio[33].gpio_I.pad_ana ;
 wire \gpio[33].gpio_I.pad_in ;
 wire \gpio[33].gpio_I.pad_oe ;
 wire \gpio[33].gpio_I.pad_out ;
 wire \gpio[34].gpio_I.pad_ana ;
 wire \gpio[34].gpio_I.pad_in ;
 wire \gpio[34].gpio_I.pad_oe ;
 wire \gpio[34].gpio_I.pad_out ;
 wire \gpio[35].gpio_I.pad_ana ;
 wire \gpio[35].gpio_I.pad_in ;
 wire \gpio[35].gpio_I.pad_oe ;
 wire \gpio[35].gpio_I.pad_out ;
 wire \gpio[36].gpio_I.pad_ana ;
 wire \gpio[36].gpio_I.pad_in ;
 wire \gpio[36].gpio_I.pad_oe ;
 wire \gpio[36].gpio_I.pad_out ;
 wire \gpio[37].gpio_I.pad_ana ;
 wire \gpio[37].gpio_I.pad_in ;
 wire \gpio[37].gpio_I.pad_oe ;
 wire \gpio[37].gpio_I.pad_out ;
 wire \gpio[38].gpio_I.pad_ana ;
 wire \gpio[38].gpio_I.pad_in ;
 wire \gpio[38].gpio_I.pad_oe ;
 wire \gpio[38].gpio_I.pad_out ;
 wire \gpio[39].gpio_I.pad_ana ;
 wire \gpio[39].gpio_I.pad_in ;
 wire \gpio[39].gpio_I.pad_oe ;
 wire \gpio[39].gpio_I.pad_out ;
 wire \gpio[3].gpio_I.pad_ana ;
 wire \gpio[3].gpio_I.pad_in ;
 wire \gpio[40].gpio_I.pad_ana ;
 wire \gpio[40].gpio_I.pad_in ;
 wire \gpio[41].gpio_I.pad_ana ;
 wire \gpio[41].gpio_I.pad_in ;
 wire \gpio[42].gpio_I.pad_ana ;
 wire \gpio[42].gpio_I.pad_in ;
 wire \gpio[43].gpio_I.pad_ana ;
 wire \gpio[43].gpio_I.pad_in ;
 wire \gpio[44].gpio_I.pad_ana ;
 wire \gpio[44].gpio_I.pad_in ;
 wire \gpio[45].gpio_I.pad_ana ;
 wire \gpio[45].gpio_I.pad_in ;
 wire \gpio[46].gpio_I.pad_ana ;
 wire \gpio[46].gpio_I.pad_in ;
 wire \gpio[47].gpio_I.pad_ana ;
 wire \gpio[47].gpio_I.pad_in ;
 wire \gpio[48].gpio_I.pad_ana ;
 wire \gpio[48].gpio_I.pad_in ;
 wire \gpio[49].gpio_I.pad_ana ;
 wire \gpio[49].gpio_I.pad_in ;
 wire \gpio[4].gpio_I.pad_ana ;
 wire \gpio[4].gpio_I.pad_in ;
 wire \gpio[52].gpio_I.pad_ana ;
 wire \gpio[52].gpio_I.pad_in ;
 wire \gpio[53].gpio_I.pad_ana ;
 wire \gpio[53].gpio_I.pad_in ;
 wire \gpio[54].gpio_I.pad_ana ;
 wire \gpio[54].gpio_I.pad_in ;
 wire \gpio[55].gpio_I.pad_ana ;
 wire \gpio[55].gpio_I.pad_in ;
 wire \gpio[58].gpio_I.pad_ana ;
 wire \gpio[58].gpio_I.pad_in ;
 wire \gpio[59].gpio_I.pad_ana ;
 wire \gpio[59].gpio_I.pad_in ;
 wire \gpio[5].gpio_I.pad_ana ;
 wire \gpio[5].gpio_I.pad_in ;
 wire \gpio[60].gpio_I.pad_ana ;
 wire \gpio[60].gpio_I.pad_in ;
 wire \gpio[61].gpio_I.pad_ana ;
 wire \gpio[61].gpio_I.pad_in ;
 wire \gpio[8].gpio_I.pad_ana ;
 wire \gpio[8].gpio_I.pad_in ;
 wire \gpio[8].gpio_I.pad_out ;
 wire \gpio[9].gpio_I.pad_ana ;
 wire \gpio[9].gpio_I.pad_in ;
 wire \gpio[9].gpio_I.pad_out ;
 wire \top_I.branch[0].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[0].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[0].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[0].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[0].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[0].check_mask.l_addr[0] ;
 wire \top_I.branch[0].check_mask.l_k_one ;
 wire \top_I.branch[0].check_mask.l_spine_iw[0] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[10] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[11] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[12] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[13] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[14] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[15] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[16] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[17] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[18] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[19] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[1] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[20] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[21] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[22] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[23] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[24] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[25] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[26] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[27] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[28] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[29] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[2] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[3] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[4] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[5] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[6] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[7] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[8] ;
 wire \top_I.branch[0].check_mask.l_spine_iw[9] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[0] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[10] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[11] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[12] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[13] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[14] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[15] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[16] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[17] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[18] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[19] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[1] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[20] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[21] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[22] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[23] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[24] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[25] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[2] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[3] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[4] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[5] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[6] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[7] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[8] ;
 wire \top_I.branch[0].check_mask.l_spine_ow[9] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[10].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[10].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[10].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[10].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[10].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[10].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[10].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[10].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[10].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[10].check_mask.l_addr[0] ;
 wire \top_I.branch[10].check_mask.l_addr[1] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[11].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[11].check_mask.l_addr[0] ;
 wire \top_I.branch[11].check_mask.l_addr[1] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[0] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[10] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[11] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[12] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[13] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[14] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[15] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[16] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[17] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[18] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[19] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[1] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[20] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[21] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[22] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[23] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[24] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[25] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[26] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[27] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[28] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[29] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[2] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[3] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[4] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[5] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[6] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[7] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[8] ;
 wire \top_I.branch[11].check_mask.l_spine_iw[9] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[0] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[10] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[11] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[12] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[13] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[14] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[15] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[16] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[17] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[18] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[19] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[1] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[20] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[21] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[22] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[23] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[24] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[25] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[2] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[3] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[4] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[5] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[6] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[7] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[8] ;
 wire \top_I.branch[11].check_mask.l_spine_ow[9] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[12].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[12].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[12].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[12].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[12].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[12].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[12].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[12].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[12].check_mask.l_addr[0] ;
 wire \top_I.branch[12].check_mask.l_addr[1] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[13].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[13].check_mask.l_addr[0] ;
 wire \top_I.branch[13].check_mask.l_addr[1] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[14].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[14].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[14].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[14].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[14].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[14].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[14].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[14].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[14].check_mask.l_addr[0] ;
 wire \top_I.branch[14].check_mask.l_addr[3] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[15].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[15].check_mask.l_addr[0] ;
 wire \top_I.branch[15].check_mask.l_addr[3] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[16].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[16].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[16].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[16].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[16].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[16].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[16].check_mask.l_addr[0] ;
 wire \top_I.branch[16].check_mask.l_addr[3] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[17].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[17].check_mask.l_addr[0] ;
 wire \top_I.branch[17].check_mask.l_addr[3] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[18].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[18].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[18].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[18].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[18].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[18].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[18].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[18].check_mask.l_addr[0] ;
 wire \top_I.branch[18].check_mask.l_addr[1] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[19].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[19].check_mask.l_addr[0] ;
 wire \top_I.branch[19].check_mask.l_addr[1] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[1].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[1].check_mask.l_addr[0] ;
 wire \top_I.branch[1].check_mask.l_k_one ;
 wire \top_I.branch[20].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[20].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[20].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[20].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[20].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[20].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[20].check_mask.l_addr[0] ;
 wire \top_I.branch[20].check_mask.l_addr[1] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[21].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[21].check_mask.l_addr[0] ;
 wire \top_I.branch[21].check_mask.l_addr[1] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[22].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[22].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[22].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[22].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[22].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[22].check_mask.l_addr[0] ;
 wire \top_I.branch[22].check_mask.l_addr[2] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[23].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[23].check_mask.l_addr[0] ;
 wire \top_I.branch[23].check_mask.l_addr[2] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[24].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[24].check_mask.l_addr[0] ;
 wire \top_I.branch[24].check_mask.l_addr[2] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[25].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[25].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[25].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[25].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[25].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[25].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[25].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[25].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[25].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[25].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[25].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[25].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[25].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[25].check_mask.l_addr[0] ;
 wire \top_I.branch[25].check_mask.l_addr[2] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[26].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[26].check_mask.l_addr[0] ;
 wire \top_I.branch[26].check_mask.l_addr[1] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[27].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[27].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[27].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[27].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[27].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[27].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[27].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[27].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[27].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[27].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[27].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[27].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[27].check_mask.l_addr[0] ;
 wire \top_I.branch[27].check_mask.l_addr[1] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[2].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[2].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[2].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[2].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[2].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[2].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[2].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[2].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[2].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[2].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[2].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[2].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[2].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[2].check_mask.l_addr[0] ;
 wire \top_I.branch[2].check_mask.l_addr[1] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[3].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[3].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[3].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[3].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[3].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[3].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[3].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[3].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[3].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[3].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[3].check_mask.l_addr[0] ;
 wire \top_I.branch[3].check_mask.l_addr[1] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[4].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[4].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[4].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[4].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[4].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[4].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[4].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[4].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[4].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[4].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[4].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[4].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[4].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[4].check_mask.l_addr[0] ;
 wire \top_I.branch[4].check_mask.l_addr[1] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[5].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[5].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[5].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[5].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[5].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[5].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[5].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[5].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[5].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[5].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[5].check_mask.l_addr[0] ;
 wire \top_I.branch[5].check_mask.l_addr[1] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[6].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[6].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[6].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[6].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[6].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[6].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[6].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[6].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[6].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[6].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[6].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[6].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[6].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[6].check_mask.l_addr[0] ;
 wire \top_I.branch[6].check_mask.l_addr[2] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[7].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[7].check_mask.l_addr[0] ;
 wire \top_I.branch[7].check_mask.l_addr[2] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[8].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[8].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[8].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[8].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[8].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[8].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[8].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[8].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[8].check_mask.l_addr[0] ;
 wire \top_I.branch[8].check_mask.l_addr[2] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[0].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[10].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[10].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[11].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[11].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[12].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[12].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[13].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[13].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[14].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[14].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[15].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[15].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[16].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[16].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[17].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[17].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[18].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[18].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[19].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[19].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[1].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[1].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[2].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[2].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[3].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[3].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[4].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[4].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[5].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[5].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[6].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[6].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[7].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[7].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[8].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[8].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.block[9].um_I.clk ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ena ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[10] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[11] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[12] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[13] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[14] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[15] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[16] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[17] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[1] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[2] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[3] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[4] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[5] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[6] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[7] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[8] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.iw[9] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.k_zero ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[0] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[10] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[11] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[12] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[13] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[14] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[15] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[16] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[17] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[18] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[19] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[1] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[20] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[21] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[22] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[23] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[2] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[3] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[4] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[5] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[6] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[7] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[8] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.ow[9] ;
 wire \top_I.branch[9].check_mask.block[9].um_I.pg_ena ;
 wire \top_I.branch[9].check_mask.l_addr[0] ;
 wire \top_I.branch[9].check_mask.l_addr[2] ;
 wire vapwr;
 wire [63:0] pad_raw;

 sg13g2_IOPadIn \gpio[0].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[0].gpio_I.pad_in ),
    .pad(pad_raw[0]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut4mA \gpio[10].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[10].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[10]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut4mA \gpio[11].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[11].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[11]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut4mA \gpio[12].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[12].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[12]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut4mA \gpio[13].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[13].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[13]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut4mA \gpio[14].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[14].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[14]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut4mA \gpio[15].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[15].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[15]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVdd \gpio[16].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[17].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[18].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[19].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[1].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[1].gpio_I.pad_in ),
    .pad(pad_raw[1]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[20].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[21].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVdd \gpio[22].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[23].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[24].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[25].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[26].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[27].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadVss \gpio[28].gpio_I.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadVdd \gpio[29].gpio_I.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[2].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[2].gpio_I.pad_in ),
    .pad(pad_raw[2]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[30].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVdd \gpio[31].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut4mA \gpio[32].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[32].gpio_I.pad_out ),
    .c2p_en(\gpio[32].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[32].gpio_I.pad_in ),
    .pad(pad_raw[32]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut4mA \gpio[33].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[33].gpio_I.pad_out ),
    .c2p_en(\gpio[33].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[33].gpio_I.pad_in ),
    .pad(pad_raw[33]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut4mA \gpio[34].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[34].gpio_I.pad_out ),
    .c2p_en(\gpio[34].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[34].gpio_I.pad_in ),
    .pad(pad_raw[34]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut4mA \gpio[35].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[35].gpio_I.pad_out ),
    .c2p_en(\gpio[35].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[35].gpio_I.pad_in ),
    .pad(pad_raw[35]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut4mA \gpio[36].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[36].gpio_I.pad_out ),
    .c2p_en(\gpio[36].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[36].gpio_I.pad_in ),
    .pad(pad_raw[36]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut4mA \gpio[37].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[37].gpio_I.pad_out ),
    .c2p_en(\gpio[37].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[37].gpio_I.pad_in ),
    .pad(pad_raw[37]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut4mA \gpio[38].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[38].gpio_I.pad_out ),
    .c2p_en(\gpio[38].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[38].gpio_I.pad_in ),
    .pad(pad_raw[38]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadInOut4mA \gpio[39].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[39].gpio_I.pad_out ),
    .c2p_en(\gpio[39].gpio_I.pad_oe ),
    .iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[39].gpio_I.pad_in ),
    .pad(pad_raw[39]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[3].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[3].gpio_I.pad_in ),
    .pad(pad_raw[3]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[40].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[40].gpio_I.pad_in ),
    .pad(pad_raw[40]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[41].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[41].gpio_I.pad_in ),
    .pad(pad_raw[41]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[42].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[42].gpio_I.pad_in ),
    .pad(pad_raw[42]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[43].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[43].gpio_I.pad_in ),
    .pad(pad_raw[43]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[44].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[44].gpio_I.pad_in ),
    .pad(pad_raw[44]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[45].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[45].gpio_I.pad_in ),
    .pad(pad_raw[45]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[46].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[46].gpio_I.pad_in ),
    .pad(pad_raw[46]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[47].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[47].gpio_I.pad_in ),
    .pad(pad_raw[47]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[48].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[48].gpio_I.pad_in ),
    .pad(pad_raw[48]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[49].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[49].gpio_I.pad_in ),
    .pad(pad_raw[49]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[4].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[4].gpio_I.pad_in ),
    .pad(pad_raw[4]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[50].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVdd \gpio[51].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[52].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[53].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[54].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[55].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[56].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVdd \gpio[57].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[58].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[59].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIn \gpio[5].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .p2c(\gpio[5].gpio_I.pad_in ),
    .pad(pad_raw[5]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[60].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[61].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadVss \gpio[62].gpio_I.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadVdd \gpio[63].gpio_I.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[6].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadIOVss \gpio[7].gpio_I.genblk1.genblk1.genblk1.pad_I  (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut4mA \gpio[8].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[8].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[8]),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_IOPadOut4mA \gpio[9].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.c2p(\gpio[9].gpio_I.pad_out ),
    .iovdd(iovdd),
    .iovss(iovss),
    .pad(pad_raw[9]),
    .vdd(vdpwr),
    .vss(vgnd));
 tt_um_chip_rom \top_I.branch[0].check_mask.block[0].um_I.block_0_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[0] }));
 tt_um_jamesrosssharp_tiny1bitam \top_I.branch[0].check_mask.block[10].um_I.block_0_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[0] }));
 tt_um_frequency_counter \top_I.branch[0].check_mask.block[12].um_I.block_0_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[0] }));
 tt_um_pid_controller \top_I.branch[0].check_mask.block[14].um_I.block_0_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[0] }));
 tt_um_rtfb_collatz \top_I.branch[0].check_mask.block[16].um_I.block_0_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[0] }));
 tt_um_wokwi_413387065339458561 \top_I.branch[0].check_mask.block[18].um_I.block_0_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[0] }));
 tt_um_factory_test \top_I.branch[0].check_mask.block[1].um_I.block_0_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[0] }));
 tt_um_tiny_ternary_tapeout_csa \top_I.branch[0].check_mask.block[2].um_I.block_0_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[0] }));
 tt_um_couchand_cora16 \top_I.branch[0].check_mask.block[4].um_I.block_0_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[0] }));
 tt_um_znah_vga_ca \top_I.branch[0].check_mask.block[6].um_I.block_0_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[0] }));
 tt_um_arandomdev_fir_engine_top \top_I.branch[0].check_mask.block[8].um_I.block_0_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[0].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[0].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[0].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[0] }));
 tt_mux \top_I.branch[0].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[0].check_mask.l_k_one ),
    .k_zero(\top_I.branch[0].check_mask.l_addr[0] ),
    .addr({\top_I.branch[0].check_mask.l_addr[0] ,
    \top_I.branch[0].check_mask.l_addr[0] ,
    \top_I.branch[0].check_mask.l_addr[0] ,
    \top_I.branch[0].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[0].check_mask.block[19].um_I.ena ,
    \top_I.branch[0].check_mask.block[18].um_I.ena ,
    \top_I.branch[0].check_mask.block[17].um_I.ena ,
    \top_I.branch[0].check_mask.block[16].um_I.ena ,
    \top_I.branch[0].check_mask.block[15].um_I.ena ,
    \top_I.branch[0].check_mask.block[14].um_I.ena ,
    \top_I.branch[0].check_mask.block[13].um_I.ena ,
    \top_I.branch[0].check_mask.block[12].um_I.ena ,
    \top_I.branch[0].check_mask.block[11].um_I.ena ,
    \top_I.branch[0].check_mask.block[10].um_I.ena ,
    \top_I.branch[0].check_mask.block[9].um_I.ena ,
    \top_I.branch[0].check_mask.block[8].um_I.ena ,
    \top_I.branch[0].check_mask.block[7].um_I.ena ,
    \top_I.branch[0].check_mask.block[6].um_I.ena ,
    \top_I.branch[0].check_mask.block[5].um_I.ena ,
    \top_I.branch[0].check_mask.block[4].um_I.ena ,
    \top_I.branch[0].check_mask.block[3].um_I.ena ,
    \top_I.branch[0].check_mask.block[2].um_I.ena ,
    \top_I.branch[0].check_mask.block[1].um_I.ena ,
    \top_I.branch[0].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[0].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[19].um_I.clk ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[18].um_I.clk ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[17].um_I.clk ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[16].um_I.clk ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[15].um_I.clk ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[14].um_I.clk ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[13].um_I.clk ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[12].um_I.clk ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[11].um_I.clk ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[10].um_I.clk ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[9].um_I.clk ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[8].um_I.clk ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[7].um_I.clk ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[6].um_I.clk ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[5].um_I.clk ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[4].um_I.clk ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[3].um_I.clk ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[2].um_I.clk ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[1].um_I.clk ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[0].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[0].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[0].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[0].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[0].check_mask.block[0].um_I.pg_ena }));
 tt_um_brukstus_tdc_with_spi \top_I.branch[10].check_mask.block[10].um_I.block_10_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[10].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[10].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[10].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[10].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[10].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[10].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[10].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[10].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[0] }));
 tt_um_iitbbs \top_I.branch[10].check_mask.block[14].um_I.block_10_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[10].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[10].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[10].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[10].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[10].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[10].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[10].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[10].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[0] }));
 tt_um_toivoh_demo_tt08 \top_I.branch[10].check_mask.block[16].um_I.block_10_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[10].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[10].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[10].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[10].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[10].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[10].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[10].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[10].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[0] }));
 tt_um_MichaelBell_canon \top_I.branch[10].check_mask.block[18].um_I.block_10_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[10].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[10].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[10].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[10].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[10].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[10].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[10].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[10].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[0] }));
 tt_um_space_invaders_game \top_I.branch[10].check_mask.block[2].um_I.block_10_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[10].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[10].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[10].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[10].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[10].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[10].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[10].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[10].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[0] }));
 tt_um_Qwendu_spi_fpu \top_I.branch[10].check_mask.block[6].um_I.block_10_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[10].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[10].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[10].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[10].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[10].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[10].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[10].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[10].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[0] }));
 tt_mux \top_I.branch[10].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[10].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[10].check_mask.l_addr[1] ),
    .addr({\top_I.branch[10].check_mask.l_addr[1] ,
    \top_I.branch[10].check_mask.l_addr[0] ,
    \top_I.branch[10].check_mask.l_addr[1] ,
    \top_I.branch[10].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[10].check_mask.block[19].um_I.ena ,
    \top_I.branch[10].check_mask.block[18].um_I.ena ,
    \top_I.branch[10].check_mask.block[17].um_I.ena ,
    \top_I.branch[10].check_mask.block[16].um_I.ena ,
    \top_I.branch[10].check_mask.block[15].um_I.ena ,
    \top_I.branch[10].check_mask.block[14].um_I.ena ,
    \top_I.branch[10].check_mask.block[13].um_I.ena ,
    \top_I.branch[10].check_mask.block[12].um_I.ena ,
    \top_I.branch[10].check_mask.block[11].um_I.ena ,
    \top_I.branch[10].check_mask.block[10].um_I.ena ,
    \top_I.branch[10].check_mask.block[9].um_I.ena ,
    \top_I.branch[10].check_mask.block[8].um_I.ena ,
    \top_I.branch[10].check_mask.block[7].um_I.ena ,
    \top_I.branch[10].check_mask.block[6].um_I.ena ,
    \top_I.branch[10].check_mask.block[5].um_I.ena ,
    \top_I.branch[10].check_mask.block[4].um_I.ena ,
    \top_I.branch[10].check_mask.block[3].um_I.ena ,
    \top_I.branch[10].check_mask.block[2].um_I.ena ,
    \top_I.branch[10].check_mask.block[1].um_I.ena ,
    \top_I.branch[10].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[10].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[19].um_I.clk ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[18].um_I.clk ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[17].um_I.clk ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[16].um_I.clk ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[15].um_I.clk ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[14].um_I.clk ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[13].um_I.clk ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[12].um_I.clk ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[11].um_I.clk ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[10].um_I.clk ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[9].um_I.clk ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[8].um_I.clk ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[7].um_I.clk ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[6].um_I.clk ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[5].um_I.clk ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[4].um_I.clk ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[3].um_I.clk ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[2].um_I.clk ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[1].um_I.clk ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[10].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[10].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[10].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[10].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[10].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[10].check_mask.block[0].um_I.pg_ena }));
 tt_um_Esteban_Oman_Mendoza_maze_2024_top \top_I.branch[11].check_mask.block[0].um_I.block_11_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[0] }));
 tt_um_juarez_jimenez \top_I.branch[11].check_mask.block[10].um_I.block_11_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[0] }));
 tt_um_control_block \top_I.branch[11].check_mask.block[11].um_I.block_11_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[0] }));
 tt_um_lif_clarencechan28 \top_I.branch[11].check_mask.block[12].um_I.block_11_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[0] }));
 tt_um_LFSR_Encrypt \top_I.branch[11].check_mask.block[13].um_I.block_11_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[0] }));
 tt_um_uart_mvm \top_I.branch[11].check_mask.block[14].um_I.block_11_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[0] }));
 tt_um_cdc_test \top_I.branch[11].check_mask.block[15].um_I.block_11_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[0] }));
 tt_um_algofoogle_tt09_ring_osc \top_I.branch[11].check_mask.block[16].um_I.block_11_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[0] }));
 tt_um_two_lif_stdp \top_I.branch[11].check_mask.block[17].um_I.block_11_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[0] }));
 tt_um_delta_liafn \top_I.branch[11].check_mask.block[18].um_I.block_11_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[0] }));
 tt_um_mikegoelzer_7segmentbyte \top_I.branch[11].check_mask.block[19].um_I.block_11_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[0] }));
 tt_um_uart_mvm_sys \top_I.branch[11].check_mask.block[1].um_I.block_11_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[0] }));
 tt_um_sebastienparadis_hamming_top \top_I.branch[11].check_mask.block[2].um_I.block_11_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[0] }));
 tt_um_MichaelBell_hd_8b10b \top_I.branch[11].check_mask.block[3].um_I.block_11_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[0] }));
 tt_um_prefix8 \top_I.branch[11].check_mask.block[4].um_I.block_11_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[0] }));
 tt_um_program_counter_top_level \top_I.branch[11].check_mask.block[5].um_I.block_11_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[0] }));
 tt_um_lif_tk \top_I.branch[11].check_mask.block[6].um_I.block_11_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[0] }));
 tt_um_murmann_group \top_I.branch[11].check_mask.block[7].um_I.block_11_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[0] }));
 tt_um_asheldon44_dsm_decimation_filter \top_I.branch[11].check_mask.block[8].um_I.block_11_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[0] }));
 tt_um_adder_accumulator_sathworld \top_I.branch[11].check_mask.block[9].um_I.block_11_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[11].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[11].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[11].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[11].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[11].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[11].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[11].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[11].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[11].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[11].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[11].check_mask.l_addr[1] ),
    .addr({\top_I.branch[11].check_mask.l_addr[1] ,
    \top_I.branch[11].check_mask.l_addr[0] ,
    \top_I.branch[11].check_mask.l_addr[1] ,
    \top_I.branch[11].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[11].check_mask.block[19].um_I.ena ,
    \top_I.branch[11].check_mask.block[18].um_I.ena ,
    \top_I.branch[11].check_mask.block[17].um_I.ena ,
    \top_I.branch[11].check_mask.block[16].um_I.ena ,
    \top_I.branch[11].check_mask.block[15].um_I.ena ,
    \top_I.branch[11].check_mask.block[14].um_I.ena ,
    \top_I.branch[11].check_mask.block[13].um_I.ena ,
    \top_I.branch[11].check_mask.block[12].um_I.ena ,
    \top_I.branch[11].check_mask.block[11].um_I.ena ,
    \top_I.branch[11].check_mask.block[10].um_I.ena ,
    \top_I.branch[11].check_mask.block[9].um_I.ena ,
    \top_I.branch[11].check_mask.block[8].um_I.ena ,
    \top_I.branch[11].check_mask.block[7].um_I.ena ,
    \top_I.branch[11].check_mask.block[6].um_I.ena ,
    \top_I.branch[11].check_mask.block[5].um_I.ena ,
    \top_I.branch[11].check_mask.block[4].um_I.ena ,
    \top_I.branch[11].check_mask.block[3].um_I.ena ,
    \top_I.branch[11].check_mask.block[2].um_I.ena ,
    \top_I.branch[11].check_mask.block[1].um_I.ena ,
    \top_I.branch[11].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[11].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[19].um_I.clk ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[18].um_I.clk ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[17].um_I.clk ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[16].um_I.clk ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[15].um_I.clk ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[14].um_I.clk ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[13].um_I.clk ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[12].um_I.clk ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[11].um_I.clk ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[10].um_I.clk ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[9].um_I.clk ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[8].um_I.clk ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[7].um_I.clk ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[6].um_I.clk ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[5].um_I.clk ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[4].um_I.clk ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[3].um_I.clk ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[2].um_I.clk ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[1].um_I.clk ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[11].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[11].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[11].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[11].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[11].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[11].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[11].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[11].check_mask.block[0].um_I.pg_ena }));
 tt_um_gfg_development_tinymandelbrot \top_I.branch[12].check_mask.block[0].um_I.block_12_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[12].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[12].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[12].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[12].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[12].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[12].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[12].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[12].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[0] }));
 tt_um_a1k0n_demo \top_I.branch[12].check_mask.block[12].um_I.block_12_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[12].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[12].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[12].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[12].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[12].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[12].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[12].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[12].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[0] }));
 tt_um_larva \top_I.branch[12].check_mask.block[18].um_I.block_12_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[12].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[12].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[12].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[12].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[12].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[12].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[12].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[12].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[0] }));
 tt_um_a1k0n_vgadonut \top_I.branch[12].check_mask.block[4].um_I.block_12_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[12].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[12].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[12].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[12].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[12].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[12].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[12].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[12].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[0] }));
 tt_um_zec_square1 \top_I.branch[12].check_mask.block[8].um_I.block_12_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[12].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[12].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[12].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[12].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[12].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[12].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[12].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[12].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[0] }));
 tt_mux \top_I.branch[12].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[12].check_mask.l_addr[1] ),
    .k_zero(\top_I.branch[12].check_mask.l_addr[0] ),
    .addr({\top_I.branch[12].check_mask.l_addr[0] ,
    \top_I.branch[12].check_mask.l_addr[1] ,
    \top_I.branch[12].check_mask.l_addr[1] ,
    \top_I.branch[12].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[12].check_mask.block[19].um_I.ena ,
    \top_I.branch[12].check_mask.block[18].um_I.ena ,
    \top_I.branch[12].check_mask.block[17].um_I.ena ,
    \top_I.branch[12].check_mask.block[16].um_I.ena ,
    \top_I.branch[12].check_mask.block[15].um_I.ena ,
    \top_I.branch[12].check_mask.block[14].um_I.ena ,
    \top_I.branch[12].check_mask.block[13].um_I.ena ,
    \top_I.branch[12].check_mask.block[12].um_I.ena ,
    \top_I.branch[12].check_mask.block[11].um_I.ena ,
    \top_I.branch[12].check_mask.block[10].um_I.ena ,
    \top_I.branch[12].check_mask.block[9].um_I.ena ,
    \top_I.branch[12].check_mask.block[8].um_I.ena ,
    \top_I.branch[12].check_mask.block[7].um_I.ena ,
    \top_I.branch[12].check_mask.block[6].um_I.ena ,
    \top_I.branch[12].check_mask.block[5].um_I.ena ,
    \top_I.branch[12].check_mask.block[4].um_I.ena ,
    \top_I.branch[12].check_mask.block[3].um_I.ena ,
    \top_I.branch[12].check_mask.block[2].um_I.ena ,
    \top_I.branch[12].check_mask.block[1].um_I.ena ,
    \top_I.branch[12].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[12].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[19].um_I.clk ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[18].um_I.clk ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[17].um_I.clk ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[16].um_I.clk ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[15].um_I.clk ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[14].um_I.clk ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[13].um_I.clk ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[12].um_I.clk ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[11].um_I.clk ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[10].um_I.clk ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[9].um_I.clk ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[8].um_I.clk ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[7].um_I.clk ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[6].um_I.clk ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[5].um_I.clk ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[4].um_I.clk ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[3].um_I.clk ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[2].um_I.clk ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[1].um_I.clk ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[12].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[12].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[12].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[12].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[12].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[12].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[12].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[12].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[12].check_mask.block[0].um_I.pg_ena }));
 tt_um_claudiotalarico_counter \top_I.branch[13].check_mask.block[0].um_I.block_13_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[0] }));
 tt_um_kashmaster_carryskip \top_I.branch[13].check_mask.block[10].um_I.block_13_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[0] }));
 tt_um_shifter \top_I.branch[13].check_mask.block[11].um_I.block_13_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[0] }));
 tt_um_wokwi_411379488132926465 \top_I.branch[13].check_mask.block[12].um_I.block_13_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[0] }));
 tt_um_lrc_stevej \top_I.branch[13].check_mask.block[13].um_I.block_13_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[0] }));
 tt_um_mroblesh \top_I.branch[13].check_mask.block[14].um_I.block_13_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[0] }));
 tt_um_tommythorn_workshop \top_I.branch[13].check_mask.block[15].um_I.block_13_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[0] }));
 tt_um_carryskip_adder9 \top_I.branch[13].check_mask.block[16].um_I.block_13_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[0] }));
 tt_um_wokwi_414120248222232577 \top_I.branch[13].check_mask.block[17].um_I.block_13_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[0] }));
 tt_um_idann \top_I.branch[13].check_mask.block[18].um_I.block_13_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[0] }));
 tt_um_tinysynth \top_I.branch[13].check_mask.block[19].um_I.block_13_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[0] }));
 tt_um_dff_mem \top_I.branch[13].check_mask.block[1].um_I.block_13_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[0] }));
 tt_um_VanceWiberg_top \top_I.branch[13].check_mask.block[2].um_I.block_13_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[0] }));
 tt_um_algofoogle_tt09_ring_osc2 \top_I.branch[13].check_mask.block[3].um_I.block_13_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[0] }));
 tt_um_ronikant_jeremykam_tinyregisters \top_I.branch[13].check_mask.block[4].um_I.block_13_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[0] }));
 tt_um_systolicLif \top_I.branch[13].check_mask.block[5].um_I.block_13_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[0] }));
 tt_um_chip4lyfe \top_I.branch[13].check_mask.block[6].um_I.block_13_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[0] }));
 tt_um_anislam \top_I.branch[13].check_mask.block[7].um_I.block_13_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[0] }));
 tt_um_array_secD7 \top_I.branch[13].check_mask.block[8].um_I.block_13_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[0] }));
 tt_um_schoeberl_test \top_I.branch[13].check_mask.block[9].um_I.block_13_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[13].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[13].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[13].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[13].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[13].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[13].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[13].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[13].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[13].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[13].check_mask.l_addr[1] ),
    .k_zero(\top_I.branch[13].check_mask.l_addr[0] ),
    .addr({\top_I.branch[13].check_mask.l_addr[0] ,
    \top_I.branch[13].check_mask.l_addr[1] ,
    \top_I.branch[13].check_mask.l_addr[1] ,
    \top_I.branch[13].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[13].check_mask.block[19].um_I.ena ,
    \top_I.branch[13].check_mask.block[18].um_I.ena ,
    \top_I.branch[13].check_mask.block[17].um_I.ena ,
    \top_I.branch[13].check_mask.block[16].um_I.ena ,
    \top_I.branch[13].check_mask.block[15].um_I.ena ,
    \top_I.branch[13].check_mask.block[14].um_I.ena ,
    \top_I.branch[13].check_mask.block[13].um_I.ena ,
    \top_I.branch[13].check_mask.block[12].um_I.ena ,
    \top_I.branch[13].check_mask.block[11].um_I.ena ,
    \top_I.branch[13].check_mask.block[10].um_I.ena ,
    \top_I.branch[13].check_mask.block[9].um_I.ena ,
    \top_I.branch[13].check_mask.block[8].um_I.ena ,
    \top_I.branch[13].check_mask.block[7].um_I.ena ,
    \top_I.branch[13].check_mask.block[6].um_I.ena ,
    \top_I.branch[13].check_mask.block[5].um_I.ena ,
    \top_I.branch[13].check_mask.block[4].um_I.ena ,
    \top_I.branch[13].check_mask.block[3].um_I.ena ,
    \top_I.branch[13].check_mask.block[2].um_I.ena ,
    \top_I.branch[13].check_mask.block[1].um_I.ena ,
    \top_I.branch[13].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[13].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[19].um_I.clk ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[18].um_I.clk ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[17].um_I.clk ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[16].um_I.clk ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[15].um_I.clk ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[14].um_I.clk ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[13].um_I.clk ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[12].um_I.clk ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[11].um_I.clk ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[10].um_I.clk ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[9].um_I.clk ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[8].um_I.clk ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[7].um_I.clk ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[6].um_I.clk ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[5].um_I.clk ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[4].um_I.clk ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[3].um_I.clk ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[2].um_I.clk ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[1].um_I.clk ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[13].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[13].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[13].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[13].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[13].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[13].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[13].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[13].check_mask.block[0].um_I.pg_ena }));
 tt_um_jayjaywong12 \top_I.branch[14].check_mask.block[10].um_I.block_14_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[14].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[14].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[14].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[14].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[14].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[14].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[14].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[14].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[0] }));
 tt_um_ddc_arghunter \top_I.branch[14].check_mask.block[14].um_I.block_14_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[14].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[14].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[14].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[14].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[14].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[14].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[14].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[14].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[0] }));
 tt_um_toivoh_demo_deluxe \top_I.branch[14].check_mask.block[18].um_I.block_14_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[14].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[14].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[14].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[14].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[14].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[14].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[14].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[14].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[0] }));
 tt_um_MichaelBell_mandelbrot \top_I.branch[14].check_mask.block[2].um_I.block_14_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[14].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[14].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[14].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[14].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[14].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[14].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[14].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[14].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[0] }));
 tt_um_silice \top_I.branch[14].check_mask.block[6].um_I.block_14_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[14].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[14].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[14].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[14].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[14].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[14].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[14].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[14].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[0] }));
 tt_mux \top_I.branch[14].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[14].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[14].check_mask.l_addr[3] ),
    .addr({\top_I.branch[14].check_mask.l_addr[3] ,
    \top_I.branch[14].check_mask.l_addr[0] ,
    \top_I.branch[14].check_mask.l_addr[0] ,
    \top_I.branch[14].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[14].check_mask.block[19].um_I.ena ,
    \top_I.branch[14].check_mask.block[18].um_I.ena ,
    \top_I.branch[14].check_mask.block[17].um_I.ena ,
    \top_I.branch[14].check_mask.block[16].um_I.ena ,
    \top_I.branch[14].check_mask.block[15].um_I.ena ,
    \top_I.branch[14].check_mask.block[14].um_I.ena ,
    \top_I.branch[14].check_mask.block[13].um_I.ena ,
    \top_I.branch[14].check_mask.block[12].um_I.ena ,
    \top_I.branch[14].check_mask.block[11].um_I.ena ,
    \top_I.branch[14].check_mask.block[10].um_I.ena ,
    \top_I.branch[14].check_mask.block[9].um_I.ena ,
    \top_I.branch[14].check_mask.block[8].um_I.ena ,
    \top_I.branch[14].check_mask.block[7].um_I.ena ,
    \top_I.branch[14].check_mask.block[6].um_I.ena ,
    \top_I.branch[14].check_mask.block[5].um_I.ena ,
    \top_I.branch[14].check_mask.block[4].um_I.ena ,
    \top_I.branch[14].check_mask.block[3].um_I.ena ,
    \top_I.branch[14].check_mask.block[2].um_I.ena ,
    \top_I.branch[14].check_mask.block[1].um_I.ena ,
    \top_I.branch[14].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[14].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[19].um_I.clk ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[18].um_I.clk ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[17].um_I.clk ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[16].um_I.clk ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[15].um_I.clk ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[14].um_I.clk ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[13].um_I.clk ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[12].um_I.clk ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[11].um_I.clk ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[10].um_I.clk ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[9].um_I.clk ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[8].um_I.clk ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[7].um_I.clk ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[6].um_I.clk ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[5].um_I.clk ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[4].um_I.clk ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[3].um_I.clk ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[2].um_I.clk ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[1].um_I.clk ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[14].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[14].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[14].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[14].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[14].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[14].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[14].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[14].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[14].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[14].check_mask.block[0].um_I.pg_ena }));
 tt_um_gmejiamtz \top_I.branch[15].check_mask.block[0].um_I.block_15_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[0] }));
 tt_um_ece298a_8_bit_cpu_top \top_I.branch[15].check_mask.block[10].um_I.block_15_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[0] }));
 tt_um_anas_7193 \top_I.branch[15].check_mask.block[11].um_I.block_15_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[0] }));
 tt_um_CarrySelect8bit \top_I.branch[15].check_mask.block[12].um_I.block_15_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[0] }));
 tt_um_flyingfish800 \top_I.branch[15].check_mask.block[13].um_I.block_15_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[0] }));
 tt_um_koggestone_adder8 \top_I.branch[15].check_mask.block[14].um_I.block_15_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[0] }));
 tt_um_project_tt09 \top_I.branch[15].check_mask.block[15].um_I.block_15_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[0] }));
 tt_um_Rapoport \top_I.branch[15].check_mask.block[16].um_I.block_15_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[0] }));
 tt_um_lifn \top_I.branch[15].check_mask.block[17].um_I.block_15_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[0] }));
 tt_um_cellular_alchemist \top_I.branch[15].check_mask.block[18].um_I.block_15_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[0] }));
 tt_um_michaelmcculloch_alu \top_I.branch[15].check_mask.block[19].um_I.block_15_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[0] }));
 tt_um_nomuwill \top_I.branch[15].check_mask.block[1].um_I.block_15_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[0] }));
 tt_um_I2C \top_I.branch[15].check_mask.block[2].um_I.block_15_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[0] }));
 tt_um_digital_clock_example \top_I.branch[15].check_mask.block[3].um_I.block_15_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[0] }));
 tt_um_perceptron_mtchun \top_I.branch[15].check_mask.block[4].um_I.block_15_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[0] }));
 tt_um_udxs \top_I.branch[15].check_mask.block[5].um_I.block_15_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[0] }));
 tt_um_histogramming \top_I.branch[15].check_mask.block[6].um_I.block_15_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[0] }));
 tt_um_matrix_mult \top_I.branch[15].check_mask.block[7].um_I.block_15_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[0] }));
 tt_um_MichaelBell_rle_vga \top_I.branch[15].check_mask.block[8].um_I.block_15_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[0] }));
 tt_um_db_MAC \top_I.branch[15].check_mask.block[9].um_I.block_15_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[15].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[15].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[15].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[15].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[15].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[15].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[15].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[15].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[15].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[15].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[15].check_mask.l_addr[3] ),
    .addr({\top_I.branch[15].check_mask.l_addr[3] ,
    \top_I.branch[15].check_mask.l_addr[0] ,
    \top_I.branch[15].check_mask.l_addr[0] ,
    \top_I.branch[15].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[15].check_mask.block[19].um_I.ena ,
    \top_I.branch[15].check_mask.block[18].um_I.ena ,
    \top_I.branch[15].check_mask.block[17].um_I.ena ,
    \top_I.branch[15].check_mask.block[16].um_I.ena ,
    \top_I.branch[15].check_mask.block[15].um_I.ena ,
    \top_I.branch[15].check_mask.block[14].um_I.ena ,
    \top_I.branch[15].check_mask.block[13].um_I.ena ,
    \top_I.branch[15].check_mask.block[12].um_I.ena ,
    \top_I.branch[15].check_mask.block[11].um_I.ena ,
    \top_I.branch[15].check_mask.block[10].um_I.ena ,
    \top_I.branch[15].check_mask.block[9].um_I.ena ,
    \top_I.branch[15].check_mask.block[8].um_I.ena ,
    \top_I.branch[15].check_mask.block[7].um_I.ena ,
    \top_I.branch[15].check_mask.block[6].um_I.ena ,
    \top_I.branch[15].check_mask.block[5].um_I.ena ,
    \top_I.branch[15].check_mask.block[4].um_I.ena ,
    \top_I.branch[15].check_mask.block[3].um_I.ena ,
    \top_I.branch[15].check_mask.block[2].um_I.ena ,
    \top_I.branch[15].check_mask.block[1].um_I.ena ,
    \top_I.branch[15].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[15].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[19].um_I.clk ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[18].um_I.clk ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[17].um_I.clk ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[16].um_I.clk ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[15].um_I.clk ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[14].um_I.clk ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[13].um_I.clk ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[12].um_I.clk ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[11].um_I.clk ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[10].um_I.clk ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[9].um_I.clk ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[8].um_I.clk ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[7].um_I.clk ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[6].um_I.clk ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[5].um_I.clk ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[4].um_I.clk ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[3].um_I.clk ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[2].um_I.clk ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[1].um_I.clk ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[15].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[15].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[15].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[15].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[15].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[15].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[15].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[15].check_mask.block[0].um_I.pg_ena }));
 tt_um_brandonramos_VGA_Pong_with_NES_Controllers \top_I.branch[16].check_mask.block[0].um_I.block_16_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[16].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[16].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[16].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[16].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[16].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[16].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[16].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[16].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[0] }));
 tt_um_bilal_trng \top_I.branch[16].check_mask.block[18].um_I.block_16_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[16].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[16].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[16].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[16].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[16].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[16].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[16].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[16].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[0] }));
 tt_um_jamesrosssharp_1bitam \top_I.branch[16].check_mask.block[6].um_I.block_16_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[16].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[16].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[16].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[16].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[16].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[16].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[16].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[16].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[0] }));
 tt_mux \top_I.branch[16].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[16].check_mask.l_addr[3] ),
    .k_zero(\top_I.branch[16].check_mask.l_addr[0] ),
    .addr({\top_I.branch[16].check_mask.l_addr[3] ,
    \top_I.branch[16].check_mask.l_addr[0] ,
    \top_I.branch[16].check_mask.l_addr[0] ,
    \top_I.branch[16].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[16].check_mask.block[19].um_I.ena ,
    \top_I.branch[16].check_mask.block[18].um_I.ena ,
    \top_I.branch[16].check_mask.block[17].um_I.ena ,
    \top_I.branch[16].check_mask.block[16].um_I.ena ,
    \top_I.branch[16].check_mask.block[15].um_I.ena ,
    \top_I.branch[16].check_mask.block[14].um_I.ena ,
    \top_I.branch[16].check_mask.block[13].um_I.ena ,
    \top_I.branch[16].check_mask.block[12].um_I.ena ,
    \top_I.branch[16].check_mask.block[11].um_I.ena ,
    \top_I.branch[16].check_mask.block[10].um_I.ena ,
    \top_I.branch[16].check_mask.block[9].um_I.ena ,
    \top_I.branch[16].check_mask.block[8].um_I.ena ,
    \top_I.branch[16].check_mask.block[7].um_I.ena ,
    \top_I.branch[16].check_mask.block[6].um_I.ena ,
    \top_I.branch[16].check_mask.block[5].um_I.ena ,
    \top_I.branch[16].check_mask.block[4].um_I.ena ,
    \top_I.branch[16].check_mask.block[3].um_I.ena ,
    \top_I.branch[16].check_mask.block[2].um_I.ena ,
    \top_I.branch[16].check_mask.block[1].um_I.ena ,
    \top_I.branch[16].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[16].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[19].um_I.clk ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[18].um_I.clk ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[17].um_I.clk ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[16].um_I.clk ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[15].um_I.clk ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[14].um_I.clk ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[13].um_I.clk ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[12].um_I.clk ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[11].um_I.clk ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[10].um_I.clk ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[9].um_I.clk ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[8].um_I.clk ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[7].um_I.clk ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[6].um_I.clk ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[5].um_I.clk ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[4].um_I.clk ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[3].um_I.clk ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[2].um_I.clk ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[1].um_I.clk ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[16].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[16].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[16].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[16].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[16].check_mask.block[0].um_I.pg_ena }));
 tt_um_kev_ma_matmult222 \top_I.branch[17].check_mask.block[0].um_I.block_17_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[0] }));
 tt_um_09eksdee \top_I.branch[17].check_mask.block[10].um_I.block_17_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[0] }));
 tt_um_urish_simon \top_I.branch[17].check_mask.block[11].um_I.block_17_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[0] }));
 tt_um_tommythorn_cgates \top_I.branch[17].check_mask.block[12].um_I.block_17_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[0] }));
 tt_um_gxrii_spi_sevenseg \top_I.branch[17].check_mask.block[13].um_I.block_17_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[0] }));
 tt_um_rejunity_sn76489 \top_I.branch[17].check_mask.block[14].um_I.block_17_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[0] }));
 tt_um_atomNPU \top_I.branch[17].check_mask.block[15].um_I.block_17_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[0] }));
 tt_um_samkho_two_channel_square_wave_generator \top_I.branch[17].check_mask.block[16].um_I.block_17_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[0] }));
 tt_um_virantha_enigma \top_I.branch[17].check_mask.block[17].um_I.block_17_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[0] }));
 tt_um_dog_BILBO \top_I.branch[17].check_mask.block[18].um_I.block_17_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[0] }));
 tt_um_synth_simple_mm \top_I.branch[17].check_mask.block[19].um_I.block_17_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[0] }));
 tt_um_tinytapeout_logo_screensaver \top_I.branch[17].check_mask.block[1].um_I.block_17_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[0] }));
 tt_um_algofoogle_tt09_ring_osc3 \top_I.branch[17].check_mask.block[2].um_I.block_17_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[0] }));
 tt_um_gamepad_pmod_demo \top_I.branch[17].check_mask.block[3].um_I.block_17_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[0] }));
 tt_um_wallento_4bit_toycpu \top_I.branch[17].check_mask.block[4].um_I.block_17_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[0] }));
 tt_um_wrapper \top_I.branch[17].check_mask.block[5].um_I.block_17_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[0] }));
 tt_um_kailinsley \top_I.branch[17].check_mask.block[6].um_I.block_17_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[0] }));
 tt_um_MAC_Accelerator_OnSachinSharma \top_I.branch[17].check_mask.block[7].um_I.block_17_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[0] }));
 tt_um_rejunity_decoder \top_I.branch[17].check_mask.block[8].um_I.block_17_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[0] }));
 tt_um_xor_encryption \top_I.branch[17].check_mask.block[9].um_I.block_17_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[17].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[17].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[17].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[17].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[17].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[17].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[17].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[17].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[17].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[17].check_mask.l_addr[3] ),
    .k_zero(\top_I.branch[17].check_mask.l_addr[0] ),
    .addr({\top_I.branch[17].check_mask.l_addr[3] ,
    \top_I.branch[17].check_mask.l_addr[0] ,
    \top_I.branch[17].check_mask.l_addr[0] ,
    \top_I.branch[17].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[17].check_mask.block[19].um_I.ena ,
    \top_I.branch[17].check_mask.block[18].um_I.ena ,
    \top_I.branch[17].check_mask.block[17].um_I.ena ,
    \top_I.branch[17].check_mask.block[16].um_I.ena ,
    \top_I.branch[17].check_mask.block[15].um_I.ena ,
    \top_I.branch[17].check_mask.block[14].um_I.ena ,
    \top_I.branch[17].check_mask.block[13].um_I.ena ,
    \top_I.branch[17].check_mask.block[12].um_I.ena ,
    \top_I.branch[17].check_mask.block[11].um_I.ena ,
    \top_I.branch[17].check_mask.block[10].um_I.ena ,
    \top_I.branch[17].check_mask.block[9].um_I.ena ,
    \top_I.branch[17].check_mask.block[8].um_I.ena ,
    \top_I.branch[17].check_mask.block[7].um_I.ena ,
    \top_I.branch[17].check_mask.block[6].um_I.ena ,
    \top_I.branch[17].check_mask.block[5].um_I.ena ,
    \top_I.branch[17].check_mask.block[4].um_I.ena ,
    \top_I.branch[17].check_mask.block[3].um_I.ena ,
    \top_I.branch[17].check_mask.block[2].um_I.ena ,
    \top_I.branch[17].check_mask.block[1].um_I.ena ,
    \top_I.branch[17].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[17].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[19].um_I.clk ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[18].um_I.clk ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[17].um_I.clk ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[16].um_I.clk ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[15].um_I.clk ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[14].um_I.clk ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[13].um_I.clk ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[12].um_I.clk ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[11].um_I.clk ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[10].um_I.clk ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[9].um_I.clk ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[8].um_I.clk ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[7].um_I.clk ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[6].um_I.clk ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[5].um_I.clk ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[4].um_I.clk ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[3].um_I.clk ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[2].um_I.clk ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[1].um_I.clk ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[17].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[17].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[17].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[17].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[17].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[17].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[17].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[17].check_mask.block[0].um_I.pg_ena }));
 tt_um_MichaelBell_tinyQV \top_I.branch[18].check_mask.block[10].um_I.block_18_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[18].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[18].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[18].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[18].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[18].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[18].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[18].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[18].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[0] }));
 tt_um_schoeberl_wildcat \top_I.branch[18].check_mask.block[16].um_I.block_18_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[18].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[18].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[18].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[18].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[18].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[18].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[18].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[18].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[0] }));
 tt_um_jmack2201 \top_I.branch[18].check_mask.block[18].um_I.block_18_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[18].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[18].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[18].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[18].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[18].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[18].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[18].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[18].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[0] }));
 tt_um_alphaonesoc \top_I.branch[18].check_mask.block[4].um_I.block_18_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[18].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[18].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[18].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[18].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[18].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[18].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[18].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[18].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[0] }));
 tt_mux \top_I.branch[18].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[18].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[18].check_mask.l_addr[1] ),
    .addr({\top_I.branch[18].check_mask.l_addr[0] ,
    \top_I.branch[18].check_mask.l_addr[1] ,
    \top_I.branch[18].check_mask.l_addr[1] ,
    \top_I.branch[18].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[18].check_mask.block[19].um_I.ena ,
    \top_I.branch[18].check_mask.block[18].um_I.ena ,
    \top_I.branch[18].check_mask.block[17].um_I.ena ,
    \top_I.branch[18].check_mask.block[16].um_I.ena ,
    \top_I.branch[18].check_mask.block[15].um_I.ena ,
    \top_I.branch[18].check_mask.block[14].um_I.ena ,
    \top_I.branch[18].check_mask.block[13].um_I.ena ,
    \top_I.branch[18].check_mask.block[12].um_I.ena ,
    \top_I.branch[18].check_mask.block[11].um_I.ena ,
    \top_I.branch[18].check_mask.block[10].um_I.ena ,
    \top_I.branch[18].check_mask.block[9].um_I.ena ,
    \top_I.branch[18].check_mask.block[8].um_I.ena ,
    \top_I.branch[18].check_mask.block[7].um_I.ena ,
    \top_I.branch[18].check_mask.block[6].um_I.ena ,
    \top_I.branch[18].check_mask.block[5].um_I.ena ,
    \top_I.branch[18].check_mask.block[4].um_I.ena ,
    \top_I.branch[18].check_mask.block[3].um_I.ena ,
    \top_I.branch[18].check_mask.block[2].um_I.ena ,
    \top_I.branch[18].check_mask.block[1].um_I.ena ,
    \top_I.branch[18].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[18].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[19].um_I.clk ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[18].um_I.clk ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[17].um_I.clk ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[16].um_I.clk ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[15].um_I.clk ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[14].um_I.clk ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[13].um_I.clk ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[12].um_I.clk ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[11].um_I.clk ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[10].um_I.clk ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[9].um_I.clk ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[8].um_I.clk ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[7].um_I.clk ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[6].um_I.clk ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[5].um_I.clk ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[4].um_I.clk ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[3].um_I.clk ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[2].um_I.clk ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[1].um_I.clk ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[18].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[18].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[18].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[18].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[18].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[18].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[18].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[18].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[18].check_mask.block[0].um_I.pg_ena }));
 tt_um_rejunity_vga_logo \top_I.branch[19].check_mask.block[0].um_I.block_19_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[0] }));
 tt_um_KoushikCSN_RISCV \top_I.branch[19].check_mask.block[10].um_I.block_19_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[0] }));
 tt_um_tappu_tobias1012 \top_I.branch[19].check_mask.block[11].um_I.block_19_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[0] }));
 tt_um_ccu_goatgate \top_I.branch[19].check_mask.block[12].um_I.block_19_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[0] }));
 tt_um_mp_lif_schor \top_I.branch[19].check_mask.block[13].um_I.block_19_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[0] }));
 tt_um_lif_ZB \top_I.branch[19].check_mask.block[14].um_I.block_19_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[0] }));
 tt_um_Strider93 \top_I.branch[19].check_mask.block[15].um_I.block_19_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[0] }));
 tt_um_z2a_rgb_mixer \top_I.branch[19].check_mask.block[16].um_I.block_19_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[0] }));
 tt_um_wokwi_422960078645704705 \top_I.branch[19].check_mask.block[17].um_I.block_19_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[0] }));
 tt_um_vga_clock \top_I.branch[19].check_mask.block[18].um_I.block_19_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[0] }));
 tt_um_keszocze_ssmcl \top_I.branch[19].check_mask.block[19].um_I.block_19_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[0] }));
 tt_um_mattvenn_spi_test \top_I.branch[19].check_mask.block[1].um_I.block_19_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[0] }));
 tt_um_liaf \top_I.branch[19].check_mask.block[2].um_I.block_19_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[0] }));
 tt_um_huffman_coder \top_I.branch[19].check_mask.block[3].um_I.block_19_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[0] }));
 tt_um_lif_network_MR \top_I.branch[19].check_mask.block[4].um_I.block_19_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[0] }));
 tt_um_multiplier_tt10 \top_I.branch[19].check_mask.block[5].um_I.block_19_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[0] }));
 tt_um_lsnn_hschweig \top_I.branch[19].check_mask.block[6].um_I.block_19_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[0] }));
 tt_um_kentrane_tinyspectrum \top_I.branch[19].check_mask.block[7].um_I.block_19_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[0] }));
 tt_um_Nishanth_RISCV \top_I.branch[19].check_mask.block[8].um_I.block_19_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[0] }));
 tt_um_i2c_regf \top_I.branch[19].check_mask.block[9].um_I.block_19_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[19].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[19].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[19].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[19].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[19].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[19].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[19].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[19].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[19].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[19].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[19].check_mask.l_addr[1] ),
    .addr({\top_I.branch[19].check_mask.l_addr[0] ,
    \top_I.branch[19].check_mask.l_addr[1] ,
    \top_I.branch[19].check_mask.l_addr[1] ,
    \top_I.branch[19].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[19].check_mask.block[19].um_I.ena ,
    \top_I.branch[19].check_mask.block[18].um_I.ena ,
    \top_I.branch[19].check_mask.block[17].um_I.ena ,
    \top_I.branch[19].check_mask.block[16].um_I.ena ,
    \top_I.branch[19].check_mask.block[15].um_I.ena ,
    \top_I.branch[19].check_mask.block[14].um_I.ena ,
    \top_I.branch[19].check_mask.block[13].um_I.ena ,
    \top_I.branch[19].check_mask.block[12].um_I.ena ,
    \top_I.branch[19].check_mask.block[11].um_I.ena ,
    \top_I.branch[19].check_mask.block[10].um_I.ena ,
    \top_I.branch[19].check_mask.block[9].um_I.ena ,
    \top_I.branch[19].check_mask.block[8].um_I.ena ,
    \top_I.branch[19].check_mask.block[7].um_I.ena ,
    \top_I.branch[19].check_mask.block[6].um_I.ena ,
    \top_I.branch[19].check_mask.block[5].um_I.ena ,
    \top_I.branch[19].check_mask.block[4].um_I.ena ,
    \top_I.branch[19].check_mask.block[3].um_I.ena ,
    \top_I.branch[19].check_mask.block[2].um_I.ena ,
    \top_I.branch[19].check_mask.block[1].um_I.ena ,
    \top_I.branch[19].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[19].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[19].um_I.clk ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[18].um_I.clk ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[17].um_I.clk ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[16].um_I.clk ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[15].um_I.clk ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[14].um_I.clk ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[13].um_I.clk ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[12].um_I.clk ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[11].um_I.clk ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[10].um_I.clk ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[9].um_I.clk ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[8].um_I.clk ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[7].um_I.clk ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[6].um_I.clk ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[5].um_I.clk ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[4].um_I.clk ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[3].um_I.clk ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[2].um_I.clk ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[1].um_I.clk ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[19].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[19].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[19].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[19].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[19].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[19].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[19].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[19].check_mask.block[0].um_I.pg_ena }));
 tt_um_ring_divider \top_I.branch[1].check_mask.block[0].um_I.block_1_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[0] }));
 tt_um_devmonk_ay8913 \top_I.branch[1].check_mask.block[11].um_I.block_1_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[0] }));
 tt_um_moody_mimosa \top_I.branch[1].check_mask.block[13].um_I.block_1_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[0] }));
 tt_um_branch_pred \top_I.branch[1].check_mask.block[15].um_I.block_1_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[0] }));
 tt_um_rejunity_ternary_dot \top_I.branch[1].check_mask.block[17].um_I.block_1_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[0] }));
 tt_um_gus16 \top_I.branch[1].check_mask.block[19].um_I.block_1_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[0] }));
 tt_um_bitty \top_I.branch[1].check_mask.block[1].um_I.block_1_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[0] }));
 tt_um_uart_bgdtanasa \top_I.branch[1].check_mask.block[3].um_I.block_1_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[0] }));
 tt_um_strau0106_simple_viii \top_I.branch[1].check_mask.block[5].um_I.block_1_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[0] }));
 tt_um_asgerwenneb \top_I.branch[1].check_mask.block[7].um_I.block_1_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[0] }));
 tt_um_toivoh_demo_tt10 \top_I.branch[1].check_mask.block[9].um_I.block_1_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[1].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[1].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[1].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[1].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[1].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[1].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[1].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[1].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[1].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[1].check_mask.l_k_one ),
    .k_zero(\top_I.branch[1].check_mask.l_addr[0] ),
    .addr({\top_I.branch[1].check_mask.l_addr[0] ,
    \top_I.branch[1].check_mask.l_addr[0] ,
    \top_I.branch[1].check_mask.l_addr[0] ,
    \top_I.branch[1].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[1].check_mask.block[19].um_I.ena ,
    \top_I.branch[1].check_mask.block[18].um_I.ena ,
    \top_I.branch[1].check_mask.block[17].um_I.ena ,
    \top_I.branch[1].check_mask.block[16].um_I.ena ,
    \top_I.branch[1].check_mask.block[15].um_I.ena ,
    \top_I.branch[1].check_mask.block[14].um_I.ena ,
    \top_I.branch[1].check_mask.block[13].um_I.ena ,
    \top_I.branch[1].check_mask.block[12].um_I.ena ,
    \top_I.branch[1].check_mask.block[11].um_I.ena ,
    \top_I.branch[1].check_mask.block[10].um_I.ena ,
    \top_I.branch[1].check_mask.block[9].um_I.ena ,
    \top_I.branch[1].check_mask.block[8].um_I.ena ,
    \top_I.branch[1].check_mask.block[7].um_I.ena ,
    \top_I.branch[1].check_mask.block[6].um_I.ena ,
    \top_I.branch[1].check_mask.block[5].um_I.ena ,
    \top_I.branch[1].check_mask.block[4].um_I.ena ,
    \top_I.branch[1].check_mask.block[3].um_I.ena ,
    \top_I.branch[1].check_mask.block[2].um_I.ena ,
    \top_I.branch[1].check_mask.block[1].um_I.ena ,
    \top_I.branch[1].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[1].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[19].um_I.clk ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[18].um_I.clk ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[17].um_I.clk ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[16].um_I.clk ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[15].um_I.clk ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[14].um_I.clk ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[13].um_I.clk ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[12].um_I.clk ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[11].um_I.clk ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[10].um_I.clk ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[9].um_I.clk ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[8].um_I.clk ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[7].um_I.clk ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[6].um_I.clk ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[5].um_I.clk ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[4].um_I.clk ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[3].um_I.clk ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[2].um_I.clk ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[1].um_I.clk ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[1].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[1].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[1].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[1].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[1].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[1].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[1].check_mask.block[0].um_I.pg_ena }));
 tt_um_urish_sic1 \top_I.branch[20].check_mask.block[18].um_I.block_20_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[20].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[20].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[20].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[20].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[20].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[20].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[20].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[20].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[0] }));
 tt_um_zoom_zoom \top_I.branch[20].check_mask.block[6].um_I.block_20_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[20].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[20].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[20].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[20].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[20].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[20].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[20].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[20].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[0] }));
 tt_mux \top_I.branch[20].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[20].check_mask.l_addr[1] ),
    .k_zero(\top_I.branch[20].check_mask.l_addr[0] ),
    .addr({\top_I.branch[20].check_mask.l_addr[1] ,
    \top_I.branch[20].check_mask.l_addr[0] ,
    \top_I.branch[20].check_mask.l_addr[1] ,
    \top_I.branch[20].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[20].check_mask.block[19].um_I.ena ,
    \top_I.branch[20].check_mask.block[18].um_I.ena ,
    \top_I.branch[20].check_mask.block[17].um_I.ena ,
    \top_I.branch[20].check_mask.block[16].um_I.ena ,
    \top_I.branch[20].check_mask.block[15].um_I.ena ,
    \top_I.branch[20].check_mask.block[14].um_I.ena ,
    \top_I.branch[20].check_mask.block[13].um_I.ena ,
    \top_I.branch[20].check_mask.block[12].um_I.ena ,
    \top_I.branch[20].check_mask.block[11].um_I.ena ,
    \top_I.branch[20].check_mask.block[10].um_I.ena ,
    \top_I.branch[20].check_mask.block[9].um_I.ena ,
    \top_I.branch[20].check_mask.block[8].um_I.ena ,
    \top_I.branch[20].check_mask.block[7].um_I.ena ,
    \top_I.branch[20].check_mask.block[6].um_I.ena ,
    \top_I.branch[20].check_mask.block[5].um_I.ena ,
    \top_I.branch[20].check_mask.block[4].um_I.ena ,
    \top_I.branch[20].check_mask.block[3].um_I.ena ,
    \top_I.branch[20].check_mask.block[2].um_I.ena ,
    \top_I.branch[20].check_mask.block[1].um_I.ena ,
    \top_I.branch[20].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[20].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[19].um_I.clk ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[18].um_I.clk ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[17].um_I.clk ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[16].um_I.clk ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[15].um_I.clk ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[14].um_I.clk ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[13].um_I.clk ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[12].um_I.clk ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[11].um_I.clk ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[10].um_I.clk ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[9].um_I.clk ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[8].um_I.clk ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[7].um_I.clk ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[6].um_I.clk ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[5].um_I.clk ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[4].um_I.clk ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[3].um_I.clk ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[2].um_I.clk ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[1].um_I.clk ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[20].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[20].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[20].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[20].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[20].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[20].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[20].check_mask.block[0].um_I.pg_ena }));
 tt_um_10_vga_crossyroad \top_I.branch[21].check_mask.block[0].um_I.block_21_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[0] }));
 tt_um_zhouzhouthezhou_adder \top_I.branch[21].check_mask.block[10].um_I.block_21_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[0] }));
 tt_um_save_buffer_hash_table \top_I.branch[21].check_mask.block[11].um_I.block_21_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[0] }));
 tt_um_torurstrom_async_lock \top_I.branch[21].check_mask.block[12].um_I.block_21_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[0] }));
 tt_um_reemashivva_fifo \top_I.branch[21].check_mask.block[13].um_I.block_21_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[0] }));
 tt_um_UartMain \top_I.branch[21].check_mask.block[14].um_I.block_21_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[0] }));
 tt_um_monishvr_fifo \top_I.branch[21].check_mask.block[15].um_I.block_21_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[0] }));
 tt_um_enjens \top_I.branch[21].check_mask.block[16].um_I.block_21_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[0] }));
 tt_um_nithishreddykvs \top_I.branch[21].check_mask.block[17].um_I.block_21_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[0] }));
 tt_um_luke_clock \top_I.branch[21].check_mask.block[18].um_I.block_21_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[0] }));
 tt_um_DaDDS \top_I.branch[21].check_mask.block[19].um_I.block_21_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[0] }));
 tt_um_ole_moller_priority_encoder_to_7_segment_decoder \top_I.branch[21].check_mask.block[1].um_I.block_21_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[0] }));
 tt_um_obriensp_jtag \top_I.branch[21].check_mask.block[2].um_I.block_21_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[0] }));
 tt_um_flummer_ltc \top_I.branch[21].check_mask.block[3].um_I.block_21_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[0] }));
 tt_um_jun1okamura_test0 \top_I.branch[21].check_mask.block[4].um_I.block_21_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[0] }));
 tt_um_tiny_shader_mole99 \top_I.branch[21].check_mask.block[5].um_I.block_21_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[0] }));
 tt_um_hpdl1414_uart_atudoroi \top_I.branch[21].check_mask.block[6].um_I.block_21_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[0] }));
 tt_um_rte_sine_synth \top_I.branch[21].check_mask.block[7].um_I.block_21_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[0] }));
 tt_um_jp_cd101_saw \top_I.branch[21].check_mask.block[8].um_I.block_21_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[0] }));
 tt_um_drum_goekce \top_I.branch[21].check_mask.block[9].um_I.block_21_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[21].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[21].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[21].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[21].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[21].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[21].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[21].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[21].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[21].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[21].check_mask.l_addr[1] ),
    .k_zero(\top_I.branch[21].check_mask.l_addr[0] ),
    .addr({\top_I.branch[21].check_mask.l_addr[1] ,
    \top_I.branch[21].check_mask.l_addr[0] ,
    \top_I.branch[21].check_mask.l_addr[1] ,
    \top_I.branch[21].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[21].check_mask.block[19].um_I.ena ,
    \top_I.branch[21].check_mask.block[18].um_I.ena ,
    \top_I.branch[21].check_mask.block[17].um_I.ena ,
    \top_I.branch[21].check_mask.block[16].um_I.ena ,
    \top_I.branch[21].check_mask.block[15].um_I.ena ,
    \top_I.branch[21].check_mask.block[14].um_I.ena ,
    \top_I.branch[21].check_mask.block[13].um_I.ena ,
    \top_I.branch[21].check_mask.block[12].um_I.ena ,
    \top_I.branch[21].check_mask.block[11].um_I.ena ,
    \top_I.branch[21].check_mask.block[10].um_I.ena ,
    \top_I.branch[21].check_mask.block[9].um_I.ena ,
    \top_I.branch[21].check_mask.block[8].um_I.ena ,
    \top_I.branch[21].check_mask.block[7].um_I.ena ,
    \top_I.branch[21].check_mask.block[6].um_I.ena ,
    \top_I.branch[21].check_mask.block[5].um_I.ena ,
    \top_I.branch[21].check_mask.block[4].um_I.ena ,
    \top_I.branch[21].check_mask.block[3].um_I.ena ,
    \top_I.branch[21].check_mask.block[2].um_I.ena ,
    \top_I.branch[21].check_mask.block[1].um_I.ena ,
    \top_I.branch[21].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[21].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[19].um_I.clk ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[18].um_I.clk ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[17].um_I.clk ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[16].um_I.clk ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[15].um_I.clk ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[14].um_I.clk ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[13].um_I.clk ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[12].um_I.clk ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[11].um_I.clk ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[10].um_I.clk ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[9].um_I.clk ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[8].um_I.clk ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[7].um_I.clk ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[6].um_I.clk ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[5].um_I.clk ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[4].um_I.clk ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[3].um_I.clk ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[2].um_I.clk ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[1].um_I.clk ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[21].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[21].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[21].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[21].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[21].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[21].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[21].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[21].check_mask.block[0].um_I.pg_ena }));
 tt_um_Coline3003_spect_top \top_I.branch[22].check_mask.block[10].um_I.block_22_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[22].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[22].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[22].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[22].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[22].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[22].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[22].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[22].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[0] }));
 tt_um_gregac_tiny_nn \top_I.branch[22].check_mask.block[18].um_I.block_22_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[22].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[22].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[22].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[22].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[22].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[22].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[22].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[22].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[0] }));
 tt_mux \top_I.branch[22].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[22].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[22].check_mask.l_addr[2] ),
    .addr({\top_I.branch[22].check_mask.l_addr[0] ,
    \top_I.branch[22].check_mask.l_addr[2] ,
    \top_I.branch[22].check_mask.l_addr[0] ,
    \top_I.branch[22].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[22].check_mask.block[19].um_I.ena ,
    \top_I.branch[22].check_mask.block[18].um_I.ena ,
    \top_I.branch[22].check_mask.block[17].um_I.ena ,
    \top_I.branch[22].check_mask.block[16].um_I.ena ,
    \top_I.branch[22].check_mask.block[15].um_I.ena ,
    \top_I.branch[22].check_mask.block[14].um_I.ena ,
    \top_I.branch[22].check_mask.block[13].um_I.ena ,
    \top_I.branch[22].check_mask.block[12].um_I.ena ,
    \top_I.branch[22].check_mask.block[11].um_I.ena ,
    \top_I.branch[22].check_mask.block[10].um_I.ena ,
    \top_I.branch[22].check_mask.block[9].um_I.ena ,
    \top_I.branch[22].check_mask.block[8].um_I.ena ,
    \top_I.branch[22].check_mask.block[7].um_I.ena ,
    \top_I.branch[22].check_mask.block[6].um_I.ena ,
    \top_I.branch[22].check_mask.block[5].um_I.ena ,
    \top_I.branch[22].check_mask.block[4].um_I.ena ,
    \top_I.branch[22].check_mask.block[3].um_I.ena ,
    \top_I.branch[22].check_mask.block[2].um_I.ena ,
    \top_I.branch[22].check_mask.block[1].um_I.ena ,
    \top_I.branch[22].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[22].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[19].um_I.clk ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[18].um_I.clk ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[17].um_I.clk ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[16].um_I.clk ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[15].um_I.clk ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[14].um_I.clk ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[13].um_I.clk ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[12].um_I.clk ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[11].um_I.clk ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[10].um_I.clk ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[9].um_I.clk ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[8].um_I.clk ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[7].um_I.clk ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[6].um_I.clk ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[5].um_I.clk ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[4].um_I.clk ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[3].um_I.clk ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[2].um_I.clk ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[1].um_I.clk ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[22].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[22].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[22].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[22].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[22].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[22].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[22].check_mask.block[0].um_I.pg_ena }));
 tt_um_sushi_demo \top_I.branch[23].check_mask.block[0].um_I.block_23_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[0] }));
 tt_um_spacewar \top_I.branch[23].check_mask.block[10].um_I.block_23_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[0] }));
 tt_um_spi_pwm_djuara \top_I.branch[23].check_mask.block[11].um_I.block_23_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[0] }));
 tt_um_log_afpm \top_I.branch[23].check_mask.block[12].um_I.block_23_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[0] }));
 tt_um_wokwi_411783629732984833 \top_I.branch[23].check_mask.block[13].um_I.block_23_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[0] }));
 tt_um_rkarl_Spiral \top_I.branch[23].check_mask.block[14].um_I.block_23_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[0] }));
 tt_um_wokwi_412635532198550529 \top_I.branch[23].check_mask.block[15].um_I.block_23_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[0] }));
 tt_um_led_jellyant \top_I.branch[23].check_mask.block[16].um_I.block_23_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[0] }));
 tt_um_wokwi_413385294512575489 \top_I.branch[23].check_mask.block[17].um_I.block_23_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[0] }));
 tt_um_project_tt10 \top_I.branch[23].check_mask.block[18].um_I.block_23_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[0] }));
 tt_um_wokwi_413387014781302785 \top_I.branch[23].check_mask.block[19].um_I.block_23_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[0] }));
 tt_um_ultra_tiny_cpu \top_I.branch[23].check_mask.block[1].um_I.block_23_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[0] }));
 tt_um_kch_cd101 \top_I.branch[23].check_mask.block[2].um_I.block_23_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[0] }));
 tt_um_aditya_patra \top_I.branch[23].check_mask.block[3].um_I.block_23_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[0] }));
 tt_um_zedulo_spitest1 \top_I.branch[23].check_mask.block[4].um_I.block_23_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[0] }));
 tt_um_4_bit_ALU \top_I.branch[23].check_mask.block[5].um_I.block_23_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[0] }));
 tt_um_daobaanh_rng \top_I.branch[23].check_mask.block[6].um_I.block_23_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[0] }));
 tt_um_htfab_checkers \top_I.branch[23].check_mask.block[7].um_I.block_23_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[0] }));
 tt_um_gcd_stephan \top_I.branch[23].check_mask.block[8].um_I.block_23_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[0] }));
 tt_um_toniklippeo \top_I.branch[23].check_mask.block[9].um_I.block_23_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[23].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[23].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[23].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[23].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[23].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[23].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[23].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[23].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[23].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[23].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[23].check_mask.l_addr[2] ),
    .addr({\top_I.branch[23].check_mask.l_addr[0] ,
    \top_I.branch[23].check_mask.l_addr[2] ,
    \top_I.branch[23].check_mask.l_addr[0] ,
    \top_I.branch[23].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[23].check_mask.block[19].um_I.ena ,
    \top_I.branch[23].check_mask.block[18].um_I.ena ,
    \top_I.branch[23].check_mask.block[17].um_I.ena ,
    \top_I.branch[23].check_mask.block[16].um_I.ena ,
    \top_I.branch[23].check_mask.block[15].um_I.ena ,
    \top_I.branch[23].check_mask.block[14].um_I.ena ,
    \top_I.branch[23].check_mask.block[13].um_I.ena ,
    \top_I.branch[23].check_mask.block[12].um_I.ena ,
    \top_I.branch[23].check_mask.block[11].um_I.ena ,
    \top_I.branch[23].check_mask.block[10].um_I.ena ,
    \top_I.branch[23].check_mask.block[9].um_I.ena ,
    \top_I.branch[23].check_mask.block[8].um_I.ena ,
    \top_I.branch[23].check_mask.block[7].um_I.ena ,
    \top_I.branch[23].check_mask.block[6].um_I.ena ,
    \top_I.branch[23].check_mask.block[5].um_I.ena ,
    \top_I.branch[23].check_mask.block[4].um_I.ena ,
    \top_I.branch[23].check_mask.block[3].um_I.ena ,
    \top_I.branch[23].check_mask.block[2].um_I.ena ,
    \top_I.branch[23].check_mask.block[1].um_I.ena ,
    \top_I.branch[23].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[23].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[19].um_I.clk ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[18].um_I.clk ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[17].um_I.clk ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[16].um_I.clk ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[15].um_I.clk ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[14].um_I.clk ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[13].um_I.clk ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[12].um_I.clk ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[11].um_I.clk ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[10].um_I.clk ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[9].um_I.clk ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[8].um_I.clk ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[7].um_I.clk ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[6].um_I.clk ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[5].um_I.clk ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[4].um_I.clk ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[3].um_I.clk ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[2].um_I.clk ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[1].um_I.clk ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[23].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[23].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[23].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[23].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[23].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[23].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[23].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[23].check_mask.block[0].um_I.pg_ena }));
 tt_um_quarren42_demoscene_top \top_I.branch[24].check_mask.block[11].um_I.block_24_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[0] }));
 tt_um_ran_DanielZhu \top_I.branch[24].check_mask.block[13].um_I.block_24_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[0] }));
 tt_um_kb2ghz_xalu \top_I.branch[24].check_mask.block[15].um_I.block_24_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[0] }));
 tt_um_mattvenn_rgb_mixer \top_I.branch[24].check_mask.block[17].um_I.block_24_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[0] }));
 tt_um_supermic_arghunter \top_I.branch[24].check_mask.block[18].um_I.block_24_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[0] }));
 tt_um_tommythorn_maxbw \top_I.branch[24].check_mask.block[19].um_I.block_24_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[0] }));
 tt_um_vga_glyph_mode \top_I.branch[24].check_mask.block[1].um_I.block_24_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[0] }));
 tt_um_find_the_damn_issue \top_I.branch[24].check_mask.block[2].um_I.block_24_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[0] }));
 tt_um_favoritohjs_scroller \top_I.branch[24].check_mask.block[3].um_I.block_24_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[0] }));
 tt_um_wokwi_407306064811090945 \top_I.branch[24].check_mask.block[5].um_I.block_24_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[0] }));
 tt_um_shuangyu_top \top_I.branch[24].check_mask.block[7].um_I.block_24_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[0] }));
 tt_um_crispy_vga \top_I.branch[24].check_mask.block[9].um_I.block_24_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[24].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[24].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[24].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[24].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[24].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[24].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[24].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[24].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[24].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[24].check_mask.l_addr[2] ),
    .k_zero(\top_I.branch[24].check_mask.l_addr[0] ),
    .addr({\top_I.branch[24].check_mask.l_addr[2] ,
    \top_I.branch[24].check_mask.l_addr[2] ,
    \top_I.branch[24].check_mask.l_addr[0] ,
    \top_I.branch[24].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[24].check_mask.block[19].um_I.ena ,
    \top_I.branch[24].check_mask.block[18].um_I.ena ,
    \top_I.branch[24].check_mask.block[17].um_I.ena ,
    \top_I.branch[24].check_mask.block[16].um_I.ena ,
    \top_I.branch[24].check_mask.block[15].um_I.ena ,
    \top_I.branch[24].check_mask.block[14].um_I.ena ,
    \top_I.branch[24].check_mask.block[13].um_I.ena ,
    \top_I.branch[24].check_mask.block[12].um_I.ena ,
    \top_I.branch[24].check_mask.block[11].um_I.ena ,
    \top_I.branch[24].check_mask.block[10].um_I.ena ,
    \top_I.branch[24].check_mask.block[9].um_I.ena ,
    \top_I.branch[24].check_mask.block[8].um_I.ena ,
    \top_I.branch[24].check_mask.block[7].um_I.ena ,
    \top_I.branch[24].check_mask.block[6].um_I.ena ,
    \top_I.branch[24].check_mask.block[5].um_I.ena ,
    \top_I.branch[24].check_mask.block[4].um_I.ena ,
    \top_I.branch[24].check_mask.block[3].um_I.ena ,
    \top_I.branch[24].check_mask.block[2].um_I.ena ,
    \top_I.branch[24].check_mask.block[1].um_I.ena ,
    \top_I.branch[24].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[24].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[19].um_I.clk ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[18].um_I.clk ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[17].um_I.clk ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[16].um_I.clk ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[15].um_I.clk ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[14].um_I.clk ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[13].um_I.clk ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[12].um_I.clk ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[11].um_I.clk ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[10].um_I.clk ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[9].um_I.clk ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[8].um_I.clk ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[7].um_I.clk ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[6].um_I.clk ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[5].um_I.clk ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[4].um_I.clk ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[3].um_I.clk ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[2].um_I.clk ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[1].um_I.clk ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[24].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[24].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[24].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[24].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[24].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[24].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[24].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[24].check_mask.block[0].um_I.pg_ena }));
 tt_um_wokwi_group_8 \top_I.branch[25].check_mask.block[0].um_I.block_25_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[25].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[25].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[25].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[25].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[25].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[25].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[25].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[25].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[0] }));
 tt_um_wokwi_group_3 \top_I.branch[25].check_mask.block[10].um_I.block_25_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[25].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[25].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[25].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[25].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[25].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[25].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[25].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[25].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[0] }));
 tt_um_wokwi_group_2 \top_I.branch[25].check_mask.block[12].um_I.block_25_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[25].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[25].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[25].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[25].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[25].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[25].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[25].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[25].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[0] }));
 tt_um_wokwi_group_1 \top_I.branch[25].check_mask.block[14].um_I.block_25_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[25].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[25].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[25].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[25].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[25].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[25].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[25].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[25].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[0] }));
 tt_um_wokwi_413387190167208961 \top_I.branch[25].check_mask.block[16].um_I.block_25_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[25].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[25].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[25].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[25].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[25].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[25].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[25].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[25].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[0] }));
 tt_um_wokwi_413387093939376129 \top_I.branch[25].check_mask.block[18].um_I.block_25_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[25].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[25].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[25].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[25].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[25].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[25].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[25].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[25].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[0] }));
 tt_um_wokwi_group_7 \top_I.branch[25].check_mask.block[2].um_I.block_25_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[25].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[25].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[25].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[25].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[25].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[25].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[25].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[25].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[0] }));
 tt_um_wokwi_group_6 \top_I.branch[25].check_mask.block[4].um_I.block_25_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[25].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[25].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[25].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[25].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[25].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[25].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[25].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[25].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[0] }));
 tt_um_wokwi_group_5 \top_I.branch[25].check_mask.block[6].um_I.block_25_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[25].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[25].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[25].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[25].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[25].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[25].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[25].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[25].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[0] }));
 tt_um_wokwi_group_4 \top_I.branch[25].check_mask.block[8].um_I.block_25_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[25].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[25].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[25].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[25].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[25].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[25].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[25].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[25].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[0] }));
 tt_mux \top_I.branch[25].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[25].check_mask.l_addr[2] ),
    .k_zero(\top_I.branch[25].check_mask.l_addr[0] ),
    .addr({\top_I.branch[25].check_mask.l_addr[2] ,
    \top_I.branch[25].check_mask.l_addr[2] ,
    \top_I.branch[25].check_mask.l_addr[0] ,
    \top_I.branch[25].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[25].check_mask.block[19].um_I.ena ,
    \top_I.branch[25].check_mask.block[18].um_I.ena ,
    \top_I.branch[25].check_mask.block[17].um_I.ena ,
    \top_I.branch[25].check_mask.block[16].um_I.ena ,
    \top_I.branch[25].check_mask.block[15].um_I.ena ,
    \top_I.branch[25].check_mask.block[14].um_I.ena ,
    \top_I.branch[25].check_mask.block[13].um_I.ena ,
    \top_I.branch[25].check_mask.block[12].um_I.ena ,
    \top_I.branch[25].check_mask.block[11].um_I.ena ,
    \top_I.branch[25].check_mask.block[10].um_I.ena ,
    \top_I.branch[25].check_mask.block[9].um_I.ena ,
    \top_I.branch[25].check_mask.block[8].um_I.ena ,
    \top_I.branch[25].check_mask.block[7].um_I.ena ,
    \top_I.branch[25].check_mask.block[6].um_I.ena ,
    \top_I.branch[25].check_mask.block[5].um_I.ena ,
    \top_I.branch[25].check_mask.block[4].um_I.ena ,
    \top_I.branch[25].check_mask.block[3].um_I.ena ,
    \top_I.branch[25].check_mask.block[2].um_I.ena ,
    \top_I.branch[25].check_mask.block[1].um_I.ena ,
    \top_I.branch[25].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[25].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[19].um_I.clk ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[18].um_I.clk ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[17].um_I.clk ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[16].um_I.clk ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[15].um_I.clk ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[14].um_I.clk ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[13].um_I.clk ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[12].um_I.clk ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[11].um_I.clk ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[10].um_I.clk ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[9].um_I.clk ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[8].um_I.clk ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[7].um_I.clk ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[6].um_I.clk ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[5].um_I.clk ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[4].um_I.clk ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[3].um_I.clk ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[2].um_I.clk ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[1].um_I.clk ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[25].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[25].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[25].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[25].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[25].check_mask.block[0].um_I.pg_ena }));
 tt_um_rejunity_atari2600 \top_I.branch[26].check_mask.block[10].um_I.block_26_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[0] }));
 tt_um_cfib_demo \top_I.branch[26].check_mask.block[11].um_I.block_26_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[0] }));
 tt_um_Richard28277 \top_I.branch[26].check_mask.block[13].um_I.block_26_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[0] }));
 tt_um_betz_morse_keyer \top_I.branch[26].check_mask.block[15].um_I.block_26_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[0] }));
 tt_um_nvious_graphics \top_I.branch[26].check_mask.block[17].um_I.block_26_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[0] }));
 tt_um_neural_navigators \top_I.branch[26].check_mask.block[18].um_I.block_26_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[0] }));
 tt_um_ezchips_calc \top_I.branch[26].check_mask.block[19].um_I.block_26_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[0] }));
 tt_um_roy1707018 \top_I.branch[26].check_mask.block[1].um_I.block_26_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[0] }));
 tt_um_sign_addsub \top_I.branch[26].check_mask.block[3].um_I.block_26_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[0] }));
 tt_um_patater_demokit \top_I.branch[26].check_mask.block[5].um_I.block_26_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[0] }));
 tt_um_demosiine_sda \top_I.branch[26].check_mask.block[7].um_I.block_26_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[0] }));
 tt_um_bytex64_munch \top_I.branch[26].check_mask.block[9].um_I.block_26_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[26].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[26].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[26].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[26].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[26].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[26].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[26].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[26].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[26].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[26].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[26].check_mask.l_addr[1] ),
    .addr({\top_I.branch[26].check_mask.l_addr[0] ,
    \top_I.branch[26].check_mask.l_addr[0] ,
    \top_I.branch[26].check_mask.l_addr[1] ,
    \top_I.branch[26].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[26].check_mask.block[19].um_I.ena ,
    \top_I.branch[26].check_mask.block[18].um_I.ena ,
    \top_I.branch[26].check_mask.block[17].um_I.ena ,
    \top_I.branch[26].check_mask.block[16].um_I.ena ,
    \top_I.branch[26].check_mask.block[15].um_I.ena ,
    \top_I.branch[26].check_mask.block[14].um_I.ena ,
    \top_I.branch[26].check_mask.block[13].um_I.ena ,
    \top_I.branch[26].check_mask.block[12].um_I.ena ,
    \top_I.branch[26].check_mask.block[11].um_I.ena ,
    \top_I.branch[26].check_mask.block[10].um_I.ena ,
    \top_I.branch[26].check_mask.block[9].um_I.ena ,
    \top_I.branch[26].check_mask.block[8].um_I.ena ,
    \top_I.branch[26].check_mask.block[7].um_I.ena ,
    \top_I.branch[26].check_mask.block[6].um_I.ena ,
    \top_I.branch[26].check_mask.block[5].um_I.ena ,
    \top_I.branch[26].check_mask.block[4].um_I.ena ,
    \top_I.branch[26].check_mask.block[3].um_I.ena ,
    \top_I.branch[26].check_mask.block[2].um_I.ena ,
    \top_I.branch[26].check_mask.block[1].um_I.ena ,
    \top_I.branch[26].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[26].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[19].um_I.clk ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[18].um_I.clk ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[17].um_I.clk ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[16].um_I.clk ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[15].um_I.clk ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[14].um_I.clk ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[13].um_I.clk ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[12].um_I.clk ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[11].um_I.clk ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[10].um_I.clk ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[9].um_I.clk ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[8].um_I.clk ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[7].um_I.clk ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[6].um_I.clk ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[5].um_I.clk ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[4].um_I.clk ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[3].um_I.clk ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[2].um_I.clk ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[1].um_I.clk ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[26].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[26].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[26].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[26].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[26].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[26].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[26].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[26].check_mask.block[0].um_I.pg_ena }));
 tt_um_wokwi_group_9 \top_I.branch[27].check_mask.block[0].um_I.block_27_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[27].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[27].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[27].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[27].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[27].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[27].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[27].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[27].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[0] }));
 tt_um_wokwi_group_13 \top_I.branch[27].check_mask.block[10].um_I.block_27_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[27].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[27].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[27].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[27].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[27].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[27].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[27].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[27].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[0] }));
 tt_um_multiplier_group_1 \top_I.branch[27].check_mask.block[12].um_I.block_27_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[27].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[27].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[27].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[27].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[27].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[27].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[27].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[27].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[0] }));
 tt_um_multiplier_group_2 \top_I.branch[27].check_mask.block[14].um_I.block_27_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[27].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[27].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[27].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[27].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[27].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[27].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[27].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[27].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[0] }));
 tt_um_multiplier_group_3 \top_I.branch[27].check_mask.block[16].um_I.block_27_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[27].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[27].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[27].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[27].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[27].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[27].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[27].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[27].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[0] }));
 tt_um_wokwi_group_10 \top_I.branch[27].check_mask.block[2].um_I.block_27_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[27].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[27].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[27].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[27].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[27].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[27].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[27].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[27].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[0] }));
 tt_um_wokwi_group_11 \top_I.branch[27].check_mask.block[4].um_I.block_27_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[27].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[27].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[27].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[27].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[27].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[27].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[27].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[27].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[0] }));
 tt_um_wokwi_group_12 \top_I.branch[27].check_mask.block[6].um_I.block_27_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[27].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[27].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[27].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[27].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[27].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[27].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[27].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[27].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[0] }));
 tt_um_tetrap_triggerer \top_I.branch[27].check_mask.block[8].um_I.block_27_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[27].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[27].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[27].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[27].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[27].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[27].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[27].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[27].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[0] }));
 tt_mux \top_I.branch[27].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[27].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[27].check_mask.l_addr[1] ),
    .addr({\top_I.branch[27].check_mask.l_addr[0] ,
    \top_I.branch[27].check_mask.l_addr[0] ,
    \top_I.branch[27].check_mask.l_addr[1] ,
    \top_I.branch[27].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[27].check_mask.block[19].um_I.ena ,
    \top_I.branch[27].check_mask.block[18].um_I.ena ,
    \top_I.branch[27].check_mask.block[17].um_I.ena ,
    \top_I.branch[27].check_mask.block[16].um_I.ena ,
    \top_I.branch[27].check_mask.block[15].um_I.ena ,
    \top_I.branch[27].check_mask.block[14].um_I.ena ,
    \top_I.branch[27].check_mask.block[13].um_I.ena ,
    \top_I.branch[27].check_mask.block[12].um_I.ena ,
    \top_I.branch[27].check_mask.block[11].um_I.ena ,
    \top_I.branch[27].check_mask.block[10].um_I.ena ,
    \top_I.branch[27].check_mask.block[9].um_I.ena ,
    \top_I.branch[27].check_mask.block[8].um_I.ena ,
    \top_I.branch[27].check_mask.block[7].um_I.ena ,
    \top_I.branch[27].check_mask.block[6].um_I.ena ,
    \top_I.branch[27].check_mask.block[5].um_I.ena ,
    \top_I.branch[27].check_mask.block[4].um_I.ena ,
    \top_I.branch[27].check_mask.block[3].um_I.ena ,
    \top_I.branch[27].check_mask.block[2].um_I.ena ,
    \top_I.branch[27].check_mask.block[1].um_I.ena ,
    \top_I.branch[27].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[27].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[19].um_I.clk ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[18].um_I.clk ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[17].um_I.clk ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[16].um_I.clk ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[15].um_I.clk ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[14].um_I.clk ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[13].um_I.clk ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[12].um_I.clk ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[11].um_I.clk ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[10].um_I.clk ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[9].um_I.clk ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[8].um_I.clk ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[7].um_I.clk ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[6].um_I.clk ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[5].um_I.clk ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[4].um_I.clk ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[3].um_I.clk ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[2].um_I.clk ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[1].um_I.clk ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[27].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[27].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[27].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[27].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[27].check_mask.block[0].um_I.pg_ena }));
 tt_um_Coline3003_top \top_I.branch[2].check_mask.block[0].um_I.block_2_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[2].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[2].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[2].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[2].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[2].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[2].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[2].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[2].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[0] }));
 tt_um_htfab_caterpillar \top_I.branch[2].check_mask.block[10].um_I.block_2_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[2].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[2].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[2].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[2].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[2].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[2].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[2].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[2].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[0] }));
 tt_um_purdue_socet_uart \top_I.branch[2].check_mask.block[12].um_I.block_2_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[2].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[2].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[2].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[2].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[2].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[2].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[2].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[2].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[0] }));
 tt_um_rejunity_ay8913 \top_I.branch[2].check_mask.block[14].um_I.block_2_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[2].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[2].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[2].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[2].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[2].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[2].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[2].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[2].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[0] }));
 tt_um_rejunity_vga_test01 \top_I.branch[2].check_mask.block[16].um_I.block_2_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[2].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[2].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[2].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[2].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[2].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[2].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[2].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[2].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[0] }));
 tt_um_warp \top_I.branch[2].check_mask.block[18].um_I.block_2_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[2].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[2].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[2].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[2].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[2].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[2].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[2].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[2].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[0] }));
 tt_um_dlmiles_dffram32x8_2r1w \top_I.branch[2].check_mask.block[2].um_I.block_2_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[2].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[2].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[2].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[2].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[2].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[2].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[2].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[2].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[0] }));
 tt_um_a1k0n_nyancat \top_I.branch[2].check_mask.block[4].um_I.block_2_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[2].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[2].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[2].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[2].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[2].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[2].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[2].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[2].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[0] }));
 tt_um_rejunity_e2m0_x_i8_matmul \top_I.branch[2].check_mask.block[6].um_I.block_2_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[2].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[2].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[2].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[2].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[2].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[2].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[2].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[2].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[0] }));
 tt_um_stochastic_integrator_tt9_CL123abc \top_I.branch[2].check_mask.block[8].um_I.block_2_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[2].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[2].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[2].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[2].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[2].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[2].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[2].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[2].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[0] }));
 tt_mux \top_I.branch[2].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[2].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[2].check_mask.l_addr[1] ),
    .addr({\top_I.branch[2].check_mask.l_addr[1] ,
    \top_I.branch[2].check_mask.l_addr[1] ,
    \top_I.branch[2].check_mask.l_addr[1] ,
    \top_I.branch[2].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[2].check_mask.block[19].um_I.ena ,
    \top_I.branch[2].check_mask.block[18].um_I.ena ,
    \top_I.branch[2].check_mask.block[17].um_I.ena ,
    \top_I.branch[2].check_mask.block[16].um_I.ena ,
    \top_I.branch[2].check_mask.block[15].um_I.ena ,
    \top_I.branch[2].check_mask.block[14].um_I.ena ,
    \top_I.branch[2].check_mask.block[13].um_I.ena ,
    \top_I.branch[2].check_mask.block[12].um_I.ena ,
    \top_I.branch[2].check_mask.block[11].um_I.ena ,
    \top_I.branch[2].check_mask.block[10].um_I.ena ,
    \top_I.branch[2].check_mask.block[9].um_I.ena ,
    \top_I.branch[2].check_mask.block[8].um_I.ena ,
    \top_I.branch[2].check_mask.block[7].um_I.ena ,
    \top_I.branch[2].check_mask.block[6].um_I.ena ,
    \top_I.branch[2].check_mask.block[5].um_I.ena ,
    \top_I.branch[2].check_mask.block[4].um_I.ena ,
    \top_I.branch[2].check_mask.block[3].um_I.ena ,
    \top_I.branch[2].check_mask.block[2].um_I.ena ,
    \top_I.branch[2].check_mask.block[1].um_I.ena ,
    \top_I.branch[2].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[2].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[19].um_I.clk ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[18].um_I.clk ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[17].um_I.clk ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[16].um_I.clk ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[15].um_I.clk ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[14].um_I.clk ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[13].um_I.clk ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[12].um_I.clk ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[11].um_I.clk ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[10].um_I.clk ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[9].um_I.clk ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[8].um_I.clk ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[7].um_I.clk ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[6].um_I.clk ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[5].um_I.clk ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[4].um_I.clk ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[3].um_I.clk ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[2].um_I.clk ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[1].um_I.clk ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[2].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[2].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[2].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[2].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[2].check_mask.block[0].um_I.pg_ena }));
 tt_um_i2c_peripheral_stevej \top_I.branch[3].check_mask.block[11].um_I.block_3_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[3].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[3].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[3].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[3].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[3].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[3].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[3].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[3].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[0] }));
 tt_um_yuri_panchul_adder_with_flow_control \top_I.branch[3].check_mask.block[13].um_I.block_3_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[3].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[3].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[3].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[3].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[3].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[3].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[3].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[3].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[0] }));
 tt_um_brailliance \top_I.branch[3].check_mask.block[15].um_I.block_3_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[3].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[3].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[3].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[3].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[3].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[3].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[3].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[3].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[0] }));
 tt_um_nyan \top_I.branch[3].check_mask.block[17].um_I.block_3_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[3].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[3].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[3].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[3].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[3].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[3].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[3].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[3].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[0] }));
 tt_um_fountaincoder_top_ad \top_I.branch[3].check_mask.block[19].um_I.block_3_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[3].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[3].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[3].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[3].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[3].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[3].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[3].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[3].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[0] }));
 tt_um_algofoogle_vga \top_I.branch[3].check_mask.block[1].um_I.block_3_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[3].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[3].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[3].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[3].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[3].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[3].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[3].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[3].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[0] }));
 tt_um_uwasic_dinogame \top_I.branch[3].check_mask.block[3].um_I.block_3_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[3].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[3].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[3].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[3].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[3].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[3].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[3].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[3].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[0] }));
 tt_um_ephrenm_tsal \top_I.branch[3].check_mask.block[5].um_I.block_3_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[3].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[3].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[3].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[3].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[3].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[3].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[3].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[3].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[0] }));
 tt_um_kapilan_alarm \top_I.branch[3].check_mask.block[7].um_I.block_3_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[3].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[3].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[3].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[3].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[3].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[3].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[3].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[3].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[0] }));
 tt_um_faramire_rotary_ring_wrapper \top_I.branch[3].check_mask.block[9].um_I.block_3_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[3].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[3].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[3].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[3].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[3].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[3].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[3].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[3].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[3].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[3].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[3].check_mask.l_addr[1] ),
    .addr({\top_I.branch[3].check_mask.l_addr[1] ,
    \top_I.branch[3].check_mask.l_addr[1] ,
    \top_I.branch[3].check_mask.l_addr[1] ,
    \top_I.branch[3].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[3].check_mask.block[19].um_I.ena ,
    \top_I.branch[3].check_mask.block[18].um_I.ena ,
    \top_I.branch[3].check_mask.block[17].um_I.ena ,
    \top_I.branch[3].check_mask.block[16].um_I.ena ,
    \top_I.branch[3].check_mask.block[15].um_I.ena ,
    \top_I.branch[3].check_mask.block[14].um_I.ena ,
    \top_I.branch[3].check_mask.block[13].um_I.ena ,
    \top_I.branch[3].check_mask.block[12].um_I.ena ,
    \top_I.branch[3].check_mask.block[11].um_I.ena ,
    \top_I.branch[3].check_mask.block[10].um_I.ena ,
    \top_I.branch[3].check_mask.block[9].um_I.ena ,
    \top_I.branch[3].check_mask.block[8].um_I.ena ,
    \top_I.branch[3].check_mask.block[7].um_I.ena ,
    \top_I.branch[3].check_mask.block[6].um_I.ena ,
    \top_I.branch[3].check_mask.block[5].um_I.ena ,
    \top_I.branch[3].check_mask.block[4].um_I.ena ,
    \top_I.branch[3].check_mask.block[3].um_I.ena ,
    \top_I.branch[3].check_mask.block[2].um_I.ena ,
    \top_I.branch[3].check_mask.block[1].um_I.ena ,
    \top_I.branch[3].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[3].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[19].um_I.clk ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[18].um_I.clk ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[17].um_I.clk ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[16].um_I.clk ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[15].um_I.clk ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[14].um_I.clk ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[13].um_I.clk ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[12].um_I.clk ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[11].um_I.clk ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[10].um_I.clk ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[9].um_I.clk ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[8].um_I.clk ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[7].um_I.clk ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[6].um_I.clk ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[5].um_I.clk ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[4].um_I.clk ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[3].um_I.clk ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[2].um_I.clk ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[1].um_I.clk ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[3].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[3].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[3].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[3].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[3].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[3].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[3].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[3].check_mask.block[0].um_I.pg_ena }));
 tt_um_hack_cpu \top_I.branch[4].check_mask.block[0].um_I.block_4_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[4].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[4].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[4].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[4].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[4].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[4].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[4].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[4].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[0] }));
 tt_um_dlfloatmac \top_I.branch[4].check_mask.block[10].um_I.block_4_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[4].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[4].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[4].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[4].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[4].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[4].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[4].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[4].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[0] }));
 tt_um_stochastic_addmultiply_CL123abc \top_I.branch[4].check_mask.block[12].um_I.block_4_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[4].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[4].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[4].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[4].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[4].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[4].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[4].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[4].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[0] }));
 tt_um_thexeno_rgbw_controller \top_I.branch[4].check_mask.block[14].um_I.block_4_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[4].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[4].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[4].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[4].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[4].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[4].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[4].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[4].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[0] }));
 tt_um_simon_cipher \top_I.branch[4].check_mask.block[16].um_I.block_4_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[4].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[4].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[4].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[4].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[4].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[4].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[4].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[4].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[0] }));
 tt_um_tt08_wirecube \top_I.branch[4].check_mask.block[18].um_I.block_4_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[4].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[4].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[4].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[4].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[4].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[4].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[4].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[4].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[0] }));
 tt_um_16_mic_beamformer_arghunter \top_I.branch[4].check_mask.block[2].um_I.block_4_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[4].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[4].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[4].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[4].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[4].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[4].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[4].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[4].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[0] }));
 tt_um_yuri_panchul_sea_battle_vga_game \top_I.branch[4].check_mask.block[4].um_I.block_4_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[4].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[4].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[4].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[4].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[4].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[4].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[4].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[4].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[0] }));
 tt_um_edwintorok \top_I.branch[4].check_mask.block[6].um_I.block_4_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[4].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[4].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[4].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[4].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[4].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[4].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[4].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[4].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[0] }));
 tt_um_yuri_panchul_schoolriscv_cpu_with_fibonacci_program \top_I.branch[4].check_mask.block[8].um_I.block_4_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[4].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[4].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[4].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[4].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[4].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[4].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[4].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[4].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[0] }));
 tt_mux \top_I.branch[4].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[4].check_mask.l_addr[1] ),
    .k_zero(\top_I.branch[4].check_mask.l_addr[0] ),
    .addr({\top_I.branch[4].check_mask.l_addr[0] ,
    \top_I.branch[4].check_mask.l_addr[0] ,
    \top_I.branch[4].check_mask.l_addr[1] ,
    \top_I.branch[4].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[4].check_mask.block[19].um_I.ena ,
    \top_I.branch[4].check_mask.block[18].um_I.ena ,
    \top_I.branch[4].check_mask.block[17].um_I.ena ,
    \top_I.branch[4].check_mask.block[16].um_I.ena ,
    \top_I.branch[4].check_mask.block[15].um_I.ena ,
    \top_I.branch[4].check_mask.block[14].um_I.ena ,
    \top_I.branch[4].check_mask.block[13].um_I.ena ,
    \top_I.branch[4].check_mask.block[12].um_I.ena ,
    \top_I.branch[4].check_mask.block[11].um_I.ena ,
    \top_I.branch[4].check_mask.block[10].um_I.ena ,
    \top_I.branch[4].check_mask.block[9].um_I.ena ,
    \top_I.branch[4].check_mask.block[8].um_I.ena ,
    \top_I.branch[4].check_mask.block[7].um_I.ena ,
    \top_I.branch[4].check_mask.block[6].um_I.ena ,
    \top_I.branch[4].check_mask.block[5].um_I.ena ,
    \top_I.branch[4].check_mask.block[4].um_I.ena ,
    \top_I.branch[4].check_mask.block[3].um_I.ena ,
    \top_I.branch[4].check_mask.block[2].um_I.ena ,
    \top_I.branch[4].check_mask.block[1].um_I.ena ,
    \top_I.branch[4].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[4].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[19].um_I.clk ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[18].um_I.clk ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[17].um_I.clk ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[16].um_I.clk ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[15].um_I.clk ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[14].um_I.clk ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[13].um_I.clk ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[12].um_I.clk ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[11].um_I.clk ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[10].um_I.clk ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[9].um_I.clk ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[8].um_I.clk ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[7].um_I.clk ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[6].um_I.clk ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[5].um_I.clk ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[4].um_I.clk ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[3].um_I.clk ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[2].um_I.clk ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[1].um_I.clk ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[4].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[4].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[4].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[4].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[4].check_mask.block[0].um_I.pg_ena }));
 tt_um_samuelm_pwm_generator \top_I.branch[5].check_mask.block[11].um_I.block_5_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[5].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[5].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[5].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[5].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[5].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[5].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[5].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[5].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[0] }));
 tt_um_dmtd_arghunter \top_I.branch[5].check_mask.block[13].um_I.block_5_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[5].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[5].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[5].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[5].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[5].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[5].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[5].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[5].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[0] }));
 tt_um_i2s_to_pwm_arghunter \top_I.branch[5].check_mask.block[15].um_I.block_5_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[5].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[5].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[5].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[5].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[5].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[5].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[5].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[5].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[0] }));
 tt_um_cejmu \top_I.branch[5].check_mask.block[17].um_I.block_5_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[5].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[5].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[5].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[5].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[5].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[5].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[5].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[5].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[0] }));
 tt_um_resfuzzy \top_I.branch[5].check_mask.block[19].um_I.block_5_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[5].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[5].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[5].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[5].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[5].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[5].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[5].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[5].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[0] }));
 tt_um_Electom_cla_4bits \top_I.branch[5].check_mask.block[1].um_I.block_5_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[5].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[5].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[5].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[5].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[5].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[5].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[5].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[5].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[0] }));
 tt_um_NicklausThompson_SkyKing \top_I.branch[5].check_mask.block[3].um_I.block_5_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[5].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[5].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[5].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[5].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[5].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[5].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[5].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[5].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[0] }));
 tt_um_top \top_I.branch[5].check_mask.block[5].um_I.block_5_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[5].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[5].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[5].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[5].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[5].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[5].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[5].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[5].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[0] }));
 tt_um_johshoff_metaballs \top_I.branch[5].check_mask.block[7].um_I.block_5_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[5].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[5].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[5].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[5].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[5].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[5].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[5].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[5].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[0] }));
 tt_um_faramire_stopwatch \top_I.branch[5].check_mask.block[9].um_I.block_5_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[5].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[5].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[5].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[5].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[5].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[5].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[5].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[5].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[5].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[5].check_mask.l_addr[1] ),
    .k_zero(\top_I.branch[5].check_mask.l_addr[0] ),
    .addr({\top_I.branch[5].check_mask.l_addr[0] ,
    \top_I.branch[5].check_mask.l_addr[0] ,
    \top_I.branch[5].check_mask.l_addr[1] ,
    \top_I.branch[5].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[5].check_mask.block[19].um_I.ena ,
    \top_I.branch[5].check_mask.block[18].um_I.ena ,
    \top_I.branch[5].check_mask.block[17].um_I.ena ,
    \top_I.branch[5].check_mask.block[16].um_I.ena ,
    \top_I.branch[5].check_mask.block[15].um_I.ena ,
    \top_I.branch[5].check_mask.block[14].um_I.ena ,
    \top_I.branch[5].check_mask.block[13].um_I.ena ,
    \top_I.branch[5].check_mask.block[12].um_I.ena ,
    \top_I.branch[5].check_mask.block[11].um_I.ena ,
    \top_I.branch[5].check_mask.block[10].um_I.ena ,
    \top_I.branch[5].check_mask.block[9].um_I.ena ,
    \top_I.branch[5].check_mask.block[8].um_I.ena ,
    \top_I.branch[5].check_mask.block[7].um_I.ena ,
    \top_I.branch[5].check_mask.block[6].um_I.ena ,
    \top_I.branch[5].check_mask.block[5].um_I.ena ,
    \top_I.branch[5].check_mask.block[4].um_I.ena ,
    \top_I.branch[5].check_mask.block[3].um_I.ena ,
    \top_I.branch[5].check_mask.block[2].um_I.ena ,
    \top_I.branch[5].check_mask.block[1].um_I.ena ,
    \top_I.branch[5].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[5].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[19].um_I.clk ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[18].um_I.clk ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[17].um_I.clk ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[16].um_I.clk ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[15].um_I.clk ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[14].um_I.clk ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[13].um_I.clk ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[12].um_I.clk ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[11].um_I.clk ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[10].um_I.clk ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[9].um_I.clk ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[8].um_I.clk ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[7].um_I.clk ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[6].um_I.clk ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[5].um_I.clk ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[4].um_I.clk ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[3].um_I.clk ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[2].um_I.clk ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[1].um_I.clk ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[5].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[5].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[5].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[5].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[5].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[5].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[5].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[5].check_mask.block[0].um_I.pg_ena }));
 tt_um_pdm_pitch_filter_arghunter \top_I.branch[6].check_mask.block[0].um_I.block_6_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[6].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[6].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[6].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[6].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[6].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[6].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[6].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[6].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[0] }));
 tt_um_dlmiles_tt08_poc_uart \top_I.branch[6].check_mask.block[10].um_I.block_6_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[6].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[6].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[6].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[6].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[6].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[6].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[6].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[6].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[0] }));
 tt_um_dendraws_donut \top_I.branch[6].check_mask.block[12].um_I.block_6_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[6].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[6].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[6].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[6].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[6].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[6].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[6].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[6].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[0] }));
 tt_um_rebeccargb_vga_pride \top_I.branch[6].check_mask.block[14].um_I.block_6_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[6].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[6].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[6].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[6].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[6].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[6].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[6].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[6].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[0] }));
 tt_um_levenshtein \top_I.branch[6].check_mask.block[16].um_I.block_6_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[6].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[6].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[6].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[6].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[6].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[6].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[6].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[6].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[0] }));
 tt_um_toivoh_pio_ram_emu_example \top_I.branch[6].check_mask.block[18].um_I.block_6_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[6].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[6].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[6].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[6].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[6].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[6].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[6].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[6].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[0] }));
 tt_um_pdm_correlator_arghunter \top_I.branch[6].check_mask.block[2].um_I.block_6_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[6].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[6].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[6].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[6].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[6].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[6].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[6].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[6].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[0] }));
 tt_um_htfab_bouncy_capsule \top_I.branch[6].check_mask.block[4].um_I.block_6_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[6].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[6].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[6].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[6].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[6].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[6].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[6].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[6].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[0] }));
 tt_um_dlmiles_poc_fskmodem_hdlctrx \top_I.branch[6].check_mask.block[6].um_I.block_6_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[6].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[6].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[6].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[6].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[6].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[6].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[6].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[6].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[0] }));
 tt_um_whynot \top_I.branch[6].check_mask.block[8].um_I.block_6_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[6].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[6].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[6].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[6].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[6].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[6].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[6].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[6].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[0] }));
 tt_mux \top_I.branch[6].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[6].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[6].check_mask.l_addr[2] ),
    .addr({\top_I.branch[6].check_mask.l_addr[2] ,
    \top_I.branch[6].check_mask.l_addr[2] ,
    \top_I.branch[6].check_mask.l_addr[0] ,
    \top_I.branch[6].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[6].check_mask.block[19].um_I.ena ,
    \top_I.branch[6].check_mask.block[18].um_I.ena ,
    \top_I.branch[6].check_mask.block[17].um_I.ena ,
    \top_I.branch[6].check_mask.block[16].um_I.ena ,
    \top_I.branch[6].check_mask.block[15].um_I.ena ,
    \top_I.branch[6].check_mask.block[14].um_I.ena ,
    \top_I.branch[6].check_mask.block[13].um_I.ena ,
    \top_I.branch[6].check_mask.block[12].um_I.ena ,
    \top_I.branch[6].check_mask.block[11].um_I.ena ,
    \top_I.branch[6].check_mask.block[10].um_I.ena ,
    \top_I.branch[6].check_mask.block[9].um_I.ena ,
    \top_I.branch[6].check_mask.block[8].um_I.ena ,
    \top_I.branch[6].check_mask.block[7].um_I.ena ,
    \top_I.branch[6].check_mask.block[6].um_I.ena ,
    \top_I.branch[6].check_mask.block[5].um_I.ena ,
    \top_I.branch[6].check_mask.block[4].um_I.ena ,
    \top_I.branch[6].check_mask.block[3].um_I.ena ,
    \top_I.branch[6].check_mask.block[2].um_I.ena ,
    \top_I.branch[6].check_mask.block[1].um_I.ena ,
    \top_I.branch[6].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[6].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[19].um_I.clk ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[18].um_I.clk ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[17].um_I.clk ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[16].um_I.clk ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[15].um_I.clk ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[14].um_I.clk ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[13].um_I.clk ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[12].um_I.clk ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[11].um_I.clk ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[10].um_I.clk ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[9].um_I.clk ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[8].um_I.clk ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[7].um_I.clk ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[6].um_I.clk ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[5].um_I.clk ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[4].um_I.clk ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[3].um_I.clk ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[2].um_I.clk ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[1].um_I.clk ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[6].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[6].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[6].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[6].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[6].check_mask.block[0].um_I.pg_ena }));
 tt_um_benpayne_ps2_decoder \top_I.branch[7].check_mask.block[10].um_I.block_7_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[0] }));
 tt_um_tmkong_rgb_mixer \top_I.branch[7].check_mask.block[11].um_I.block_7_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[0] }));
 tt_um_meriac_play_tune \top_I.branch[7].check_mask.block[12].um_I.block_7_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[0] }));
 tt_um_led_matrix_ayla_lin \top_I.branch[7].check_mask.block[13].um_I.block_7_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[0] }));
 tt_um_daosvik_aesinvsbox \top_I.branch[7].check_mask.block[14].um_I.block_7_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[0] }));
 tt_um_rebeccargb_tt09ball_screensaver \top_I.branch[7].check_mask.block[15].um_I.block_7_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[0] }));
 tt_um_cattuto_sr_latch \top_I.branch[7].check_mask.block[16].um_I.block_7_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[0] }));
 tt_um_rebeccargb_colorbars \top_I.branch[7].check_mask.block[17].um_I.block_7_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[0] }));
 tt_um_emmyxu_obstacle_detection \top_I.branch[7].check_mask.block[18].um_I.block_7_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[0] }));
 tt_um_rebeccargb_hardware_utf8 \top_I.branch[7].check_mask.block[19].um_I.block_7_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[0] }));
 tt_um_vga_cbtest \top_I.branch[7].check_mask.block[1].um_I.block_7_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[0] }));
 tt_um_dpmunit \top_I.branch[7].check_mask.block[3].um_I.block_7_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[0] }));
 tt_um_mac \top_I.branch[7].check_mask.block[4].um_I.block_7_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[0] }));
 tt_um_clock_divider_arghunter \top_I.branch[7].check_mask.block[5].um_I.block_7_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[0] }));
 tt_um_dpmu \top_I.branch[7].check_mask.block[6].um_I.block_7_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[0] }));
 tt_um_emilian_muxpga \top_I.branch[7].check_mask.block[7].um_I.block_7_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[0] }));
 tt_um_JAC_EE_segdecode \top_I.branch[7].check_mask.block[8].um_I.block_7_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[0] }));
 tt_um_pyamnihc_dummy_counter \top_I.branch[7].check_mask.block[9].um_I.block_7_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[7].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[7].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[7].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[7].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[7].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[7].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[7].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[7].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[7].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[7].check_mask.l_addr[0] ),
    .k_zero(\top_I.branch[7].check_mask.l_addr[2] ),
    .addr({\top_I.branch[7].check_mask.l_addr[2] ,
    \top_I.branch[7].check_mask.l_addr[2] ,
    \top_I.branch[7].check_mask.l_addr[0] ,
    \top_I.branch[7].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[7].check_mask.block[19].um_I.ena ,
    \top_I.branch[7].check_mask.block[18].um_I.ena ,
    \top_I.branch[7].check_mask.block[17].um_I.ena ,
    \top_I.branch[7].check_mask.block[16].um_I.ena ,
    \top_I.branch[7].check_mask.block[15].um_I.ena ,
    \top_I.branch[7].check_mask.block[14].um_I.ena ,
    \top_I.branch[7].check_mask.block[13].um_I.ena ,
    \top_I.branch[7].check_mask.block[12].um_I.ena ,
    \top_I.branch[7].check_mask.block[11].um_I.ena ,
    \top_I.branch[7].check_mask.block[10].um_I.ena ,
    \top_I.branch[7].check_mask.block[9].um_I.ena ,
    \top_I.branch[7].check_mask.block[8].um_I.ena ,
    \top_I.branch[7].check_mask.block[7].um_I.ena ,
    \top_I.branch[7].check_mask.block[6].um_I.ena ,
    \top_I.branch[7].check_mask.block[5].um_I.ena ,
    \top_I.branch[7].check_mask.block[4].um_I.ena ,
    \top_I.branch[7].check_mask.block[3].um_I.ena ,
    \top_I.branch[7].check_mask.block[2].um_I.ena ,
    \top_I.branch[7].check_mask.block[1].um_I.ena ,
    \top_I.branch[7].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[7].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[19].um_I.clk ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[18].um_I.clk ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[17].um_I.clk ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[16].um_I.clk ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[15].um_I.clk ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[14].um_I.clk ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[13].um_I.clk ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[12].um_I.clk ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[11].um_I.clk ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[10].um_I.clk ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[9].um_I.clk ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[8].um_I.clk ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[7].um_I.clk ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[6].um_I.clk ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[5].um_I.clk ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[4].um_I.clk ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[3].um_I.clk ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[2].um_I.clk ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[1].um_I.clk ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[7].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[7].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[7].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[7].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[7].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[7].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[7].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[7].check_mask.block[0].um_I.pg_ena }));
 tt_um_underserved \top_I.branch[8].check_mask.block[10].um_I.block_8_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[8].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[8].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[8].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[8].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[8].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[8].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[8].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[8].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[0] }));
 tt_um_devinatkin_basys3_uart \top_I.branch[8].check_mask.block[14].um_I.block_8_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[8].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[8].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[8].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[8].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[8].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[8].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[8].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[8].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[0] }));
 tt_um_wokwi_413386991502909441 \top_I.branch[8].check_mask.block[18].um_I.block_8_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[8].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[8].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[8].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[8].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[8].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[8].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[8].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[8].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[0] }));
 tt_um_2048_vga_game \top_I.branch[8].check_mask.block[2].um_I.block_8_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[8].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[8].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[8].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[8].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[8].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[8].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[8].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[8].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[0] }));
 tt_um_rejunity_z80 \top_I.branch[8].check_mask.block[6].um_I.block_8_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[8].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[8].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[8].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[8].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[8].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[8].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[8].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[8].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[0] }));
 tt_mux \top_I.branch[8].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[8].check_mask.l_addr[2] ),
    .k_zero(\top_I.branch[8].check_mask.l_addr[0] ),
    .addr({\top_I.branch[8].check_mask.l_addr[0] ,
    \top_I.branch[8].check_mask.l_addr[2] ,
    \top_I.branch[8].check_mask.l_addr[0] ,
    \top_I.branch[8].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[8].check_mask.block[19].um_I.ena ,
    \top_I.branch[8].check_mask.block[18].um_I.ena ,
    \top_I.branch[8].check_mask.block[17].um_I.ena ,
    \top_I.branch[8].check_mask.block[16].um_I.ena ,
    \top_I.branch[8].check_mask.block[15].um_I.ena ,
    \top_I.branch[8].check_mask.block[14].um_I.ena ,
    \top_I.branch[8].check_mask.block[13].um_I.ena ,
    \top_I.branch[8].check_mask.block[12].um_I.ena ,
    \top_I.branch[8].check_mask.block[11].um_I.ena ,
    \top_I.branch[8].check_mask.block[10].um_I.ena ,
    \top_I.branch[8].check_mask.block[9].um_I.ena ,
    \top_I.branch[8].check_mask.block[8].um_I.ena ,
    \top_I.branch[8].check_mask.block[7].um_I.ena ,
    \top_I.branch[8].check_mask.block[6].um_I.ena ,
    \top_I.branch[8].check_mask.block[5].um_I.ena ,
    \top_I.branch[8].check_mask.block[4].um_I.ena ,
    \top_I.branch[8].check_mask.block[3].um_I.ena ,
    \top_I.branch[8].check_mask.block[2].um_I.ena ,
    \top_I.branch[8].check_mask.block[1].um_I.ena ,
    \top_I.branch[8].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[8].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[19].um_I.clk ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[18].um_I.clk ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[17].um_I.clk ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[16].um_I.clk ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[15].um_I.clk ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[14].um_I.clk ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[13].um_I.clk ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[12].um_I.clk ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[11].um_I.clk ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[10].um_I.clk ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[9].um_I.clk ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[8].um_I.clk ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[7].um_I.clk ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[6].um_I.clk ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[5].um_I.clk ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[4].um_I.clk ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[3].um_I.clk ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[2].um_I.clk ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[1].um_I.clk ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[8].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[8].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[8].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[8].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[8].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[8].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[8].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero ,
    \top_I.branch[8].check_mask.block[0].um_I.k_zero }),
    .um_pg_ena({\top_I.branch[8].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[8].check_mask.block[0].um_I.pg_ena }));
 tt_um_senolgulgonul \top_I.branch[9].check_mask.block[0].um_I.block_9_0.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[0].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[0].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[0] }));
 tt_um_tobimckellar_top \top_I.branch[9].check_mask.block[10].um_I.block_9_10.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[10].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[10].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[10].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[0] }));
 tt_um_alif \top_I.branch[9].check_mask.block[11].um_I.block_9_11.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[11].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[11].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[0] }));
 tt_um_rebeccargb_intercal_alu \top_I.branch[9].check_mask.block[12].um_I.block_9_12.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[12].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[12].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[12].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[0] }));
 tt_um_lif1 \top_I.branch[9].check_mask.block[13].um_I.block_9_13.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[13].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[13].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[0] }));
 tt_um_rebeccargb_universal_decoder \top_I.branch[9].check_mask.block[14].um_I.block_9_14.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[14].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[14].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[0] }));
 tt_um_instrumented_ring_oscillator \top_I.branch[9].check_mask.block[15].um_I.block_9_15.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[15].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[15].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[0] }));
 tt_um_rebeccargb_vga_timing_experiments \top_I.branch[9].check_mask.block[16].um_I.block_9_16.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[16].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[16].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[16].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[0] }));
 tt_um_lfsr_stevej \top_I.branch[9].check_mask.block[17].um_I.block_9_17.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[17].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[17].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[17].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[0] }));
 tt_um_rebeccargb_styler \top_I.branch[9].check_mask.block[18].um_I.block_9_18.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[18].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[18].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[18].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[0] }));
 tt_um_pwm_top \top_I.branch[9].check_mask.block[19].um_I.block_9_19.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[19].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[19].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[19].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[0] }));
 tt_um_hybrid_adder \top_I.branch[9].check_mask.block[1].um_I.block_9_1.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[1].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[1].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[0] }));
 tt_um_alf19185_ALU \top_I.branch[9].check_mask.block[2].um_I.block_9_2.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[2].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[2].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[0] }));
 tt_um_CLA8 \top_I.branch[9].check_mask.block[3].um_I.block_9_3.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[3].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[3].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[0] }));
 tt_um_my_elevator \top_I.branch[9].check_mask.block[4].um_I.block_9_4.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[4].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[4].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[0] }));
 tt_um_riscv_mini \top_I.branch[9].check_mask.block[5].um_I.block_9_5.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[5].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[5].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[0] }));
 tt_um_led_cipher \top_I.branch[9].check_mask.block[6].um_I.block_9_6.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[6].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[6].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[0] }));
 tt_um_carryskip_adder8 \top_I.branch[9].check_mask.block[7].um_I.block_9_7.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[7].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[7].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[0] }));
 tt_um_JesusMinguillon_freqSweep \top_I.branch[9].check_mask.block[8].um_I.block_9_8.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[8].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[8].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[0] }));
 tt_um_tiny_ternary_tapeout \top_I.branch[9].check_mask.block[9].um_I.block_9_9.tt_um_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .clk(\top_I.branch[9].check_mask.block[9].um_I.clk ),
    .ena(\top_I.branch[9].check_mask.block[9].um_I.ena ),
    .rst_n(\top_I.branch[9].check_mask.block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[9].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[9].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[9].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[9].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[9].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[9].check_mask.mux_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .k_one(\top_I.branch[9].check_mask.l_addr[2] ),
    .k_zero(\top_I.branch[9].check_mask.l_addr[0] ),
    .addr({\top_I.branch[9].check_mask.l_addr[0] ,
    \top_I.branch[9].check_mask.l_addr[2] ,
    \top_I.branch[9].check_mask.l_addr[0] ,
    \top_I.branch[9].check_mask.l_addr[0] }),
    .spine_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }),
    .um_ena({\top_I.branch[9].check_mask.block[19].um_I.ena ,
    \top_I.branch[9].check_mask.block[18].um_I.ena ,
    \top_I.branch[9].check_mask.block[17].um_I.ena ,
    \top_I.branch[9].check_mask.block[16].um_I.ena ,
    \top_I.branch[9].check_mask.block[15].um_I.ena ,
    \top_I.branch[9].check_mask.block[14].um_I.ena ,
    \top_I.branch[9].check_mask.block[13].um_I.ena ,
    \top_I.branch[9].check_mask.block[12].um_I.ena ,
    \top_I.branch[9].check_mask.block[11].um_I.ena ,
    \top_I.branch[9].check_mask.block[10].um_I.ena ,
    \top_I.branch[9].check_mask.block[9].um_I.ena ,
    \top_I.branch[9].check_mask.block[8].um_I.ena ,
    \top_I.branch[9].check_mask.block[7].um_I.ena ,
    \top_I.branch[9].check_mask.block[6].um_I.ena ,
    \top_I.branch[9].check_mask.block[5].um_I.ena ,
    \top_I.branch[9].check_mask.block[4].um_I.ena ,
    \top_I.branch[9].check_mask.block[3].um_I.ena ,
    \top_I.branch[9].check_mask.block[2].um_I.ena ,
    \top_I.branch[9].check_mask.block[1].um_I.ena ,
    \top_I.branch[9].check_mask.block[0].um_I.ena }),
    .um_iw({\top_I.branch[9].check_mask.block[19].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[19].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[19].um_I.clk ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[18].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[18].um_I.clk ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[17].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[17].um_I.clk ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[16].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[16].um_I.clk ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[15].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[15].um_I.clk ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[14].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[14].um_I.clk ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[13].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[13].um_I.clk ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[12].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[12].um_I.clk ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[11].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[11].um_I.clk ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[10].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[10].um_I.clk ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[9].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[9].um_I.clk ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[8].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[8].um_I.clk ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[7].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[7].um_I.clk ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[6].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[6].um_I.clk ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[5].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[5].um_I.clk ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[4].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[4].um_I.clk ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[3].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[3].um_I.clk ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[2].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[2].um_I.clk ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[1].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[1].um_I.clk ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[17] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[16] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[15] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[14] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[13] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[12] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[11] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[10] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[9] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[8] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[7] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[6] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[5] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[4] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[3] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[2] ,
    \top_I.branch[9].check_mask.block[0].um_I.iw[1] ,
    \top_I.branch[9].check_mask.block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[9].check_mask.block[19].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[18].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[17].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[16].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[15].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[14].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[13].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[12].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[11].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[10].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[9].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[8].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[7].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[6].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[5].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[4].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[3].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[2].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[1].um_I.k_zero ,
    \top_I.branch[9].check_mask.block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[9].check_mask.block[19].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[19].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[18].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[17].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[16].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[15].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[14].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[13].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[12].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[11].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[10].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[9].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[8].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[7].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[6].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[5].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[4].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[3].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[2].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[1].um_I.ow[0] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[23] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[22] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[21] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[20] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[19] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[18] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[17] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[16] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[15] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[14] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[13] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[12] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[11] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[10] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[9] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[8] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[7] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[6] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[5] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[4] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[3] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[2] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[1] ,
    \top_I.branch[9].check_mask.block[0].um_I.ow[0] }),
    .um_pg_ena({\top_I.branch[9].check_mask.block[19].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[18].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[17].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[16].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[15].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[14].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[13].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[12].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[11].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[10].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[9].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[8].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[7].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[6].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[5].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[4].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[3].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[2].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[1].um_I.pg_ena ,
    \top_I.branch[9].check_mask.block[0].um_I.pg_ena }));
 tt_ctrl \top_I.ctrl_I  (.VGND(vgnd),
    .VPWR(vdpwr),
    .ctrl_ena(\gpio[0].gpio_I.pad_in ),
    .ctrl_sel_inc(\gpio[1].gpio_I.pad_in ),
    .ctrl_sel_rst_n(\gpio[2].gpio_I.pad_in ),
    .k_one(\gpio[0].gpio_I.pad_oe ),
    .k_zero(\gpio[18].gpio_I.pad_oe ),
    .pad_ui_in({\gpio[47].gpio_I.pad_in ,
    \gpio[46].gpio_I.pad_in ,
    \gpio[45].gpio_I.pad_in ,
    \gpio[44].gpio_I.pad_in ,
    \gpio[43].gpio_I.pad_in ,
    \gpio[42].gpio_I.pad_in ,
    \gpio[41].gpio_I.pad_in ,
    \gpio[40].gpio_I.pad_in ,
    \gpio[48].gpio_I.pad_in ,
    \gpio[49].gpio_I.pad_in }),
    .pad_uio_in({\gpio[39].gpio_I.pad_in ,
    \gpio[38].gpio_I.pad_in ,
    \gpio[37].gpio_I.pad_in ,
    \gpio[36].gpio_I.pad_in ,
    \gpio[35].gpio_I.pad_in ,
    \gpio[34].gpio_I.pad_in ,
    \gpio[33].gpio_I.pad_in ,
    \gpio[32].gpio_I.pad_in }),
    .pad_uio_oex({\gpio[39].gpio_I.pad_oe ,
    \gpio[38].gpio_I.pad_oe ,
    \gpio[37].gpio_I.pad_oe ,
    \gpio[36].gpio_I.pad_oe ,
    \gpio[35].gpio_I.pad_oe ,
    \gpio[34].gpio_I.pad_oe ,
    \gpio[33].gpio_I.pad_oe ,
    \gpio[32].gpio_I.pad_oe }),
    .pad_uio_out({\gpio[39].gpio_I.pad_out ,
    \gpio[38].gpio_I.pad_out ,
    \gpio[37].gpio_I.pad_out ,
    \gpio[36].gpio_I.pad_out ,
    \gpio[35].gpio_I.pad_out ,
    \gpio[34].gpio_I.pad_out ,
    \gpio[33].gpio_I.pad_out ,
    \gpio[32].gpio_I.pad_out }),
    .pad_uo_out({\gpio[15].gpio_I.pad_out ,
    \gpio[14].gpio_I.pad_out ,
    \gpio[13].gpio_I.pad_out ,
    \gpio[12].gpio_I.pad_out ,
    \gpio[11].gpio_I.pad_out ,
    \gpio[10].gpio_I.pad_out ,
    \gpio[9].gpio_I.pad_out ,
    \gpio[8].gpio_I.pad_out }),
    .spine_bot_iw({\top_I.branch[0].check_mask.l_spine_iw[29] ,
    \top_I.branch[0].check_mask.l_spine_iw[28] ,
    \top_I.branch[0].check_mask.l_spine_iw[27] ,
    \top_I.branch[0].check_mask.l_spine_iw[26] ,
    \top_I.branch[0].check_mask.l_spine_iw[25] ,
    \top_I.branch[0].check_mask.l_spine_iw[24] ,
    \top_I.branch[0].check_mask.l_spine_iw[23] ,
    \top_I.branch[0].check_mask.l_spine_iw[22] ,
    \top_I.branch[0].check_mask.l_spine_iw[21] ,
    \top_I.branch[0].check_mask.l_spine_iw[20] ,
    \top_I.branch[0].check_mask.l_spine_iw[19] ,
    \top_I.branch[0].check_mask.l_spine_iw[18] ,
    \top_I.branch[0].check_mask.l_spine_iw[17] ,
    \top_I.branch[0].check_mask.l_spine_iw[16] ,
    \top_I.branch[0].check_mask.l_spine_iw[15] ,
    \top_I.branch[0].check_mask.l_spine_iw[14] ,
    \top_I.branch[0].check_mask.l_spine_iw[13] ,
    \top_I.branch[0].check_mask.l_spine_iw[12] ,
    \top_I.branch[0].check_mask.l_spine_iw[11] ,
    \top_I.branch[0].check_mask.l_spine_iw[10] ,
    \top_I.branch[0].check_mask.l_spine_iw[9] ,
    \top_I.branch[0].check_mask.l_spine_iw[8] ,
    \top_I.branch[0].check_mask.l_spine_iw[7] ,
    \top_I.branch[0].check_mask.l_spine_iw[6] ,
    \top_I.branch[0].check_mask.l_spine_iw[5] ,
    \top_I.branch[0].check_mask.l_spine_iw[4] ,
    \top_I.branch[0].check_mask.l_spine_iw[3] ,
    \top_I.branch[0].check_mask.l_spine_iw[2] ,
    \top_I.branch[0].check_mask.l_spine_iw[1] ,
    \top_I.branch[0].check_mask.l_spine_iw[0] }),
    .spine_bot_ow({\top_I.branch[0].check_mask.l_spine_ow[25] ,
    \top_I.branch[0].check_mask.l_spine_ow[24] ,
    \top_I.branch[0].check_mask.l_spine_ow[23] ,
    \top_I.branch[0].check_mask.l_spine_ow[22] ,
    \top_I.branch[0].check_mask.l_spine_ow[21] ,
    \top_I.branch[0].check_mask.l_spine_ow[20] ,
    \top_I.branch[0].check_mask.l_spine_ow[19] ,
    \top_I.branch[0].check_mask.l_spine_ow[18] ,
    \top_I.branch[0].check_mask.l_spine_ow[17] ,
    \top_I.branch[0].check_mask.l_spine_ow[16] ,
    \top_I.branch[0].check_mask.l_spine_ow[15] ,
    \top_I.branch[0].check_mask.l_spine_ow[14] ,
    \top_I.branch[0].check_mask.l_spine_ow[13] ,
    \top_I.branch[0].check_mask.l_spine_ow[12] ,
    \top_I.branch[0].check_mask.l_spine_ow[11] ,
    \top_I.branch[0].check_mask.l_spine_ow[10] ,
    \top_I.branch[0].check_mask.l_spine_ow[9] ,
    \top_I.branch[0].check_mask.l_spine_ow[8] ,
    \top_I.branch[0].check_mask.l_spine_ow[7] ,
    \top_I.branch[0].check_mask.l_spine_ow[6] ,
    \top_I.branch[0].check_mask.l_spine_ow[5] ,
    \top_I.branch[0].check_mask.l_spine_ow[4] ,
    \top_I.branch[0].check_mask.l_spine_ow[3] ,
    \top_I.branch[0].check_mask.l_spine_ow[2] ,
    \top_I.branch[0].check_mask.l_spine_ow[1] ,
    \top_I.branch[0].check_mask.l_spine_ow[0] }),
    .spine_top_iw({\top_I.branch[11].check_mask.l_spine_iw[29] ,
    \top_I.branch[11].check_mask.l_spine_iw[28] ,
    \top_I.branch[11].check_mask.l_spine_iw[27] ,
    \top_I.branch[11].check_mask.l_spine_iw[26] ,
    \top_I.branch[11].check_mask.l_spine_iw[25] ,
    \top_I.branch[11].check_mask.l_spine_iw[24] ,
    \top_I.branch[11].check_mask.l_spine_iw[23] ,
    \top_I.branch[11].check_mask.l_spine_iw[22] ,
    \top_I.branch[11].check_mask.l_spine_iw[21] ,
    \top_I.branch[11].check_mask.l_spine_iw[20] ,
    \top_I.branch[11].check_mask.l_spine_iw[19] ,
    \top_I.branch[11].check_mask.l_spine_iw[18] ,
    \top_I.branch[11].check_mask.l_spine_iw[17] ,
    \top_I.branch[11].check_mask.l_spine_iw[16] ,
    \top_I.branch[11].check_mask.l_spine_iw[15] ,
    \top_I.branch[11].check_mask.l_spine_iw[14] ,
    \top_I.branch[11].check_mask.l_spine_iw[13] ,
    \top_I.branch[11].check_mask.l_spine_iw[12] ,
    \top_I.branch[11].check_mask.l_spine_iw[11] ,
    \top_I.branch[11].check_mask.l_spine_iw[10] ,
    \top_I.branch[11].check_mask.l_spine_iw[9] ,
    \top_I.branch[11].check_mask.l_spine_iw[8] ,
    \top_I.branch[11].check_mask.l_spine_iw[7] ,
    \top_I.branch[11].check_mask.l_spine_iw[6] ,
    \top_I.branch[11].check_mask.l_spine_iw[5] ,
    \top_I.branch[11].check_mask.l_spine_iw[4] ,
    \top_I.branch[11].check_mask.l_spine_iw[3] ,
    \top_I.branch[11].check_mask.l_spine_iw[2] ,
    \top_I.branch[11].check_mask.l_spine_iw[1] ,
    \top_I.branch[11].check_mask.l_spine_iw[0] }),
    .spine_top_ow({\top_I.branch[11].check_mask.l_spine_ow[25] ,
    \top_I.branch[11].check_mask.l_spine_ow[24] ,
    \top_I.branch[11].check_mask.l_spine_ow[23] ,
    \top_I.branch[11].check_mask.l_spine_ow[22] ,
    \top_I.branch[11].check_mask.l_spine_ow[21] ,
    \top_I.branch[11].check_mask.l_spine_ow[20] ,
    \top_I.branch[11].check_mask.l_spine_ow[19] ,
    \top_I.branch[11].check_mask.l_spine_ow[18] ,
    \top_I.branch[11].check_mask.l_spine_ow[17] ,
    \top_I.branch[11].check_mask.l_spine_ow[16] ,
    \top_I.branch[11].check_mask.l_spine_ow[15] ,
    \top_I.branch[11].check_mask.l_spine_ow[14] ,
    \top_I.branch[11].check_mask.l_spine_ow[13] ,
    \top_I.branch[11].check_mask.l_spine_ow[12] ,
    \top_I.branch[11].check_mask.l_spine_ow[11] ,
    \top_I.branch[11].check_mask.l_spine_ow[10] ,
    \top_I.branch[11].check_mask.l_spine_ow[9] ,
    \top_I.branch[11].check_mask.l_spine_ow[8] ,
    \top_I.branch[11].check_mask.l_spine_ow[7] ,
    \top_I.branch[11].check_mask.l_spine_ow[6] ,
    \top_I.branch[11].check_mask.l_spine_ow[5] ,
    \top_I.branch[11].check_mask.l_spine_ow[4] ,
    \top_I.branch[11].check_mask.l_spine_ow[3] ,
    \top_I.branch[11].check_mask.l_spine_ow[2] ,
    \top_I.branch[11].check_mask.l_spine_ow[1] ,
    \top_I.branch[11].check_mask.l_spine_ow[0] }));
 sg13g2_Corner IO_CORNER_NORTH_WEST_INST (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Corner IO_CORNER_NORTH_EAST_INST (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Corner IO_CORNER_SOUTH_WEST_INST (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Corner IO_CORNER_SOUTH_EAST_INST (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_0_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_0_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_NORTH_0_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_0_120 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_1_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_1_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_1_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_1_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_1_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_1_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_2_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_2_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_2_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_2_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_2_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_2_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_3_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_3_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_3_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_3_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_3_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_3_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_4_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_4_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_4_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_4_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_4_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_4_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_5_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_5_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_5_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_5_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_5_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_5_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_6_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_6_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_6_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_6_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_6_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_6_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_7_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_7_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_7_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_7_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_7_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_7_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_8_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_8_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_8_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_8_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_8_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_8_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_9_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_9_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_9_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_9_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_9_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_9_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_10_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_10_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_10_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_10_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_10_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_10_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_11_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_11_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_11_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_11_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_11_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_11_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_12_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_12_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_12_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_12_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_12_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_12_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_13_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_13_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_13_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_13_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_13_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_13_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_14_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_NORTH_14_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_NORTH_14_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_NORTH_14_120 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_0_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_0_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_SOUTH_0_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_0_120 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_1_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_1_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_1_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_1_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_1_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_1_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_2_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_2_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_2_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_2_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_2_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_2_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_3_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_3_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_3_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_3_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_3_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_3_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_4_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_4_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_4_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_4_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_4_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_4_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_5_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_5_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_5_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_5_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_5_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_5_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_6_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_6_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_6_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_6_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_6_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_6_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_7_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_7_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_7_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_7_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_7_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_7_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_8_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_8_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_8_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_8_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_8_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_8_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_9_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_9_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_9_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_9_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_9_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_9_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_10_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_10_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_10_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_10_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_10_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_10_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_11_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_11_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_11_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_11_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_11_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_11_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_12_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_12_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_12_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_12_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_12_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_12_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_13_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_13_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_13_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_13_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_13_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_13_250 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_14_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_14_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_SOUTH_14_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_14_120 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_0_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_0_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_0_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler200 IO_FILL_IO_WEST_0_120 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_1_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_1_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_1_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_1_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_1_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_1_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_1_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_2_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_2_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_2_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_2_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_2_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_2_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_2_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_3_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_3_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_3_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_3_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_3_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_3_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_3_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_4_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_4_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_4_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_4_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_4_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_4_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_4_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_5_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_5_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_5_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_5_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_5_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_5_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_5_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_6_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_6_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_6_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_6_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_6_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_6_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_6_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_7_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_7_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_7_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_7_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_7_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_7_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_7_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_8_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_8_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_8_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_8_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_8_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_8_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_8_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_9_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_9_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_9_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_9_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_9_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_9_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_9_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_10_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_10_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_10_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_10_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_10_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_10_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_10_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_11_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_11_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_11_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_11_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_11_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_11_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_11_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_12_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_12_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_12_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_12_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_12_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_12_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_12_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_13_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_13_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_13_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_13_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_13_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_13_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_13_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_14_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_14_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_14_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_14_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_14_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_14_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_14_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_15_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_15_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_15_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_15_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_15_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_15_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_15_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_16_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_16_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_16_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_16_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_16_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_16_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_16_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_17_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_17_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_17_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_17_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_17_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_17_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_WEST_17_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_18_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_WEST_18_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_WEST_18_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_WEST_18_120 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler1000 IO_FILL_IO_WEST_18_130 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_0_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_0_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_0_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler200 IO_FILL_IO_EAST_0_120 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_1_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_1_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_1_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_1_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_1_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_1_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_1_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_2_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_2_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_2_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_2_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_2_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_2_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_2_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_3_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_3_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_3_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_3_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_3_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_3_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_3_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_4_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_4_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_4_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_4_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_4_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_4_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_4_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_5_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_5_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_5_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_5_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_5_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_5_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_5_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_6_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_6_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_6_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_6_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_6_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_6_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_6_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_7_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_7_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_7_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_7_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_7_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_7_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_7_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_8_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_8_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_8_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_8_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_8_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_8_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_8_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_9_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_9_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_9_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_9_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_9_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_9_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_9_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_10_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_10_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_10_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_10_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_10_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_10_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_10_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_11_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_11_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_11_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_11_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_11_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_11_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_11_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_12_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_12_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_12_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_12_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_12_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_12_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_12_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_13_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_13_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_13_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_13_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_13_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_13_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_13_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_14_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_14_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_14_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_14_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_14_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_14_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_14_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_15_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_15_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_15_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_15_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_15_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_15_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_15_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_16_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_16_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_16_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_16_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_16_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_16_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_16_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_17_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_17_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_17_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_17_150 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_17_200 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_17_220 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler400 IO_FILL_IO_EAST_17_240 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_18_0 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler10000 IO_FILL_IO_EAST_18_50 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler4000 IO_FILL_IO_EAST_18_100 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler2000 IO_FILL_IO_EAST_18_120 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 sg13g2_Filler1000 IO_FILL_IO_EAST_18_130 (.iovdd(iovdd),
    .iovss(iovss),
    .vdd(vdpwr),
    .vss(vgnd));
 bondpad_70x70 \IO_BOND_gpio[0].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[0]));
 bondpad_70x70 \IO_BOND_gpio[10].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[10]));
 bondpad_70x70 \IO_BOND_gpio[11].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[11]));
 bondpad_70x70 \IO_BOND_gpio[12].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[12]));
 bondpad_70x70 \IO_BOND_gpio[13].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[13]));
 bondpad_70x70 \IO_BOND_gpio[14].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[14]));
 bondpad_70x70 \IO_BOND_gpio[15].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[15]));
 bondpad_70x70 \IO_BOND_gpio[16].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(iovdd));
 bondpad_70x70 \IO_BOND_gpio[17].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[18].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[19].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[1].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[1]));
 bondpad_70x70 \IO_BOND_gpio[20].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[21].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[22].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(iovdd));
 bondpad_70x70 \IO_BOND_gpio[23].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[24].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[25].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[26].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[27].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[28].gpio_I.genblk1.pad_I  (.pad(vgnd));
 bondpad_70x70 \IO_BOND_gpio[29].gpio_I.genblk1.genblk1.pad_I  (.pad(vdpwr));
 bondpad_70x70 \IO_BOND_gpio[2].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[2]));
 bondpad_70x70 \IO_BOND_gpio[30].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[31].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(iovdd));
 bondpad_70x70 \IO_BOND_gpio[32].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[32]));
 bondpad_70x70 \IO_BOND_gpio[33].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[33]));
 bondpad_70x70 \IO_BOND_gpio[34].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[34]));
 bondpad_70x70 \IO_BOND_gpio[35].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[35]));
 bondpad_70x70 \IO_BOND_gpio[36].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[36]));
 bondpad_70x70 \IO_BOND_gpio[37].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[37]));
 bondpad_70x70 \IO_BOND_gpio[38].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[38]));
 bondpad_70x70 \IO_BOND_gpio[39].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[39]));
 bondpad_70x70 \IO_BOND_gpio[3].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[3]));
 bondpad_70x70 \IO_BOND_gpio[40].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[40]));
 bondpad_70x70 \IO_BOND_gpio[41].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[41]));
 bondpad_70x70 \IO_BOND_gpio[42].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[42]));
 bondpad_70x70 \IO_BOND_gpio[43].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[43]));
 bondpad_70x70 \IO_BOND_gpio[44].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[44]));
 bondpad_70x70 \IO_BOND_gpio[45].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[45]));
 bondpad_70x70 \IO_BOND_gpio[46].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[46]));
 bondpad_70x70 \IO_BOND_gpio[47].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[47]));
 bondpad_70x70 \IO_BOND_gpio[48].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[48]));
 bondpad_70x70 \IO_BOND_gpio[49].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[49]));
 bondpad_70x70 \IO_BOND_gpio[4].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[4]));
 bondpad_70x70 \IO_BOND_gpio[50].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[51].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(iovdd));
 bondpad_70x70 \IO_BOND_gpio[52].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[53].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[54].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[55].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[56].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[57].gpio_I.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(iovdd));
 bondpad_70x70 \IO_BOND_gpio[58].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[59].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[5].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[5]));
 bondpad_70x70 \IO_BOND_gpio[60].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[61].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[62].gpio_I.genblk1.pad_I  (.pad(vgnd));
 bondpad_70x70 \IO_BOND_gpio[63].gpio_I.genblk1.genblk1.pad_I  (.pad(vdpwr));
 bondpad_70x70 \IO_BOND_gpio[6].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[7].gpio_I.genblk1.genblk1.genblk1.pad_I  (.pad(iovss));
 bondpad_70x70 \IO_BOND_gpio[8].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[8]));
 bondpad_70x70 \IO_BOND_gpio[9].gpio_I.genblk1.genblk1.genblk1.genblk1.genblk1.genblk1.pad_I  (.pad(pad_raw[9]));
endmodule
